------------------------------------------------------------------
--  File        : fir_filter.vhd
--  Description : FIR filter
------------------------------------------------------------------
-- Filter Specifications:
--
-- Sample Rate     : 25 MHz
-- Response        : Lowpass
-- Specification   : Fp,Fst,Ap,Ast
-- Stopband Atten. : 40 dB
-- Stopband Edge   : 300 kHz
-- Passband Edge   : 200 kHz
-- Passband Ripple : 0.01 dB
----------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fir_filter is
  port (
    I_CLK : in std_logic;
    I_RST : in std_logic;
    I_FILTER : in std_logic_vector(31 downto 0);
    O_FILTER : out std_logic_vector(44 downto 0)
  );
end entity fir_filter;

architecture rtl of fir_filter is

  -- Local Functions
  -- Type Definitions
  TYPE delay_pipeline_type IS ARRAY (NATURAL range <>) OF signed(31 DOWNTO 0); -- sfix32_En31
  -- Constants
  CONSTANT coeff1                         : signed(7 DOWNTO 0) := to_signed(13, 8); -- sfix8_En12
  CONSTANT coeff2                         : signed(7 DOWNTO 0) := to_signed(-8, 8); -- sfix8_En12
  CONSTANT coeff3                         : signed(7 DOWNTO 0) := to_signed(-6, 8); -- sfix8_En12
  CONSTANT coeff4                         : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff5                         : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff6                         : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff7                         : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff8                         : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff9                         : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff10                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff11                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff12                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff13                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff14                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff15                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff16                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff17                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff18                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff19                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff20                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff21                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff22                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff23                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff24                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff25                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff26                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff27                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff28                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff29                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff30                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff31                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff32                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff33                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff34                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff35                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff36                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff37                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff38                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff39                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff40                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff41                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff42                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff43                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff44                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff45                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff46                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff47                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff48                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff49                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff50                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff51                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff52                        : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff53                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff54                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff55                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff56                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff57                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff58                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff59                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff60                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff61                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff62                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff63                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff64                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff65                        : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff66                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff67                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff68                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff69                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff70                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff71                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff72                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff73                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff74                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff75                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff76                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff77                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff78                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff79                        : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff80                        : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff81                        : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff82                        : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff83                        : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff84                        : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff85                        : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff86                        : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff87                        : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff88                        : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff89                        : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff90                        : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff91                        : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff92                        : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff93                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff94                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff95                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff96                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff97                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff98                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff99                        : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff100                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff101                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff102                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff103                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff104                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff105                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff106                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff107                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff108                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff109                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff110                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff111                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff112                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff113                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff114                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff115                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff116                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff117                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff118                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff119                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff120                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff121                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff122                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff123                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff124                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff125                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff126                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff127                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff128                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff129                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff130                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff131                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff132                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff133                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff134                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff135                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff136                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff137                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff138                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff139                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff140                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff141                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff142                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff143                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff144                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff145                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff146                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff147                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff148                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff149                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff150                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff151                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff152                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff153                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff154                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff155                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff156                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff157                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff158                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff159                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff160                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff161                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff162                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff163                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff164                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff165                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff166                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff167                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff168                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff169                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff170                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff171                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff172                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff173                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff174                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff175                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff176                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff177                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff178                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff179                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff180                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff181                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff182                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff183                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff184                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff185                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff186                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff187                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff188                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff189                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff190                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff191                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff192                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff193                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff194                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff195                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff196                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff197                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff198                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff199                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff200                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff201                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff202                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff203                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff204                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff205                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff206                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff207                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff208                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff209                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff210                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff211                       : signed(7 DOWNTO 0) := to_signed(4, 8); -- sfix8_En12
  CONSTANT coeff212                       : signed(7 DOWNTO 0) := to_signed(4, 8); -- sfix8_En12
  CONSTANT coeff213                       : signed(7 DOWNTO 0) := to_signed(5, 8); -- sfix8_En12
  CONSTANT coeff214                       : signed(7 DOWNTO 0) := to_signed(5, 8); -- sfix8_En12
  CONSTANT coeff215                       : signed(7 DOWNTO 0) := to_signed(6, 8); -- sfix8_En12
  CONSTANT coeff216                       : signed(7 DOWNTO 0) := to_signed(6, 8); -- sfix8_En12
  CONSTANT coeff217                       : signed(7 DOWNTO 0) := to_signed(6, 8); -- sfix8_En12
  CONSTANT coeff218                       : signed(7 DOWNTO 0) := to_signed(7, 8); -- sfix8_En12
  CONSTANT coeff219                       : signed(7 DOWNTO 0) := to_signed(7, 8); -- sfix8_En12
  CONSTANT coeff220                       : signed(7 DOWNTO 0) := to_signed(7, 8); -- sfix8_En12
  CONSTANT coeff221                       : signed(7 DOWNTO 0) := to_signed(8, 8); -- sfix8_En12
  CONSTANT coeff222                       : signed(7 DOWNTO 0) := to_signed(8, 8); -- sfix8_En12
  CONSTANT coeff223                       : signed(7 DOWNTO 0) := to_signed(8, 8); -- sfix8_En12
  CONSTANT coeff224                       : signed(7 DOWNTO 0) := to_signed(8, 8); -- sfix8_En12
  CONSTANT coeff225                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff226                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff227                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff228                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff229                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff230                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff231                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff232                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff233                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff234                       : signed(7 DOWNTO 0) := to_signed(8, 8); -- sfix8_En12
  CONSTANT coeff235                       : signed(7 DOWNTO 0) := to_signed(8, 8); -- sfix8_En12
  CONSTANT coeff236                       : signed(7 DOWNTO 0) := to_signed(8, 8); -- sfix8_En12
  CONSTANT coeff237                       : signed(7 DOWNTO 0) := to_signed(8, 8); -- sfix8_En12
  CONSTANT coeff238                       : signed(7 DOWNTO 0) := to_signed(7, 8); -- sfix8_En12
  CONSTANT coeff239                       : signed(7 DOWNTO 0) := to_signed(7, 8); -- sfix8_En12
  CONSTANT coeff240                       : signed(7 DOWNTO 0) := to_signed(7, 8); -- sfix8_En12
  CONSTANT coeff241                       : signed(7 DOWNTO 0) := to_signed(6, 8); -- sfix8_En12
  CONSTANT coeff242                       : signed(7 DOWNTO 0) := to_signed(6, 8); -- sfix8_En12
  CONSTANT coeff243                       : signed(7 DOWNTO 0) := to_signed(5, 8); -- sfix8_En12
  CONSTANT coeff244                       : signed(7 DOWNTO 0) := to_signed(5, 8); -- sfix8_En12
  CONSTANT coeff245                       : signed(7 DOWNTO 0) := to_signed(4, 8); -- sfix8_En12
  CONSTANT coeff246                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff247                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff248                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff249                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff250                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff251                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff252                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff253                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff254                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff255                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff256                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff257                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff258                       : signed(7 DOWNTO 0) := to_signed(-6, 8); -- sfix8_En12
  CONSTANT coeff259                       : signed(7 DOWNTO 0) := to_signed(-7, 8); -- sfix8_En12
  CONSTANT coeff260                       : signed(7 DOWNTO 0) := to_signed(-8, 8); -- sfix8_En12
  CONSTANT coeff261                       : signed(7 DOWNTO 0) := to_signed(-8, 8); -- sfix8_En12
  CONSTANT coeff262                       : signed(7 DOWNTO 0) := to_signed(-9, 8); -- sfix8_En12
  CONSTANT coeff263                       : signed(7 DOWNTO 0) := to_signed(-10, 8); -- sfix8_En12
  CONSTANT coeff264                       : signed(7 DOWNTO 0) := to_signed(-11, 8); -- sfix8_En12
  CONSTANT coeff265                       : signed(7 DOWNTO 0) := to_signed(-11, 8); -- sfix8_En12
  CONSTANT coeff266                       : signed(7 DOWNTO 0) := to_signed(-12, 8); -- sfix8_En12
  CONSTANT coeff267                       : signed(7 DOWNTO 0) := to_signed(-13, 8); -- sfix8_En12
  CONSTANT coeff268                       : signed(7 DOWNTO 0) := to_signed(-14, 8); -- sfix8_En12
  CONSTANT coeff269                       : signed(7 DOWNTO 0) := to_signed(-14, 8); -- sfix8_En12
  CONSTANT coeff270                       : signed(7 DOWNTO 0) := to_signed(-15, 8); -- sfix8_En12
  CONSTANT coeff271                       : signed(7 DOWNTO 0) := to_signed(-15, 8); -- sfix8_En12
  CONSTANT coeff272                       : signed(7 DOWNTO 0) := to_signed(-16, 8); -- sfix8_En12
  CONSTANT coeff273                       : signed(7 DOWNTO 0) := to_signed(-16, 8); -- sfix8_En12
  CONSTANT coeff274                       : signed(7 DOWNTO 0) := to_signed(-16, 8); -- sfix8_En12
  CONSTANT coeff275                       : signed(7 DOWNTO 0) := to_signed(-17, 8); -- sfix8_En12
  CONSTANT coeff276                       : signed(7 DOWNTO 0) := to_signed(-17, 8); -- sfix8_En12
  CONSTANT coeff277                       : signed(7 DOWNTO 0) := to_signed(-17, 8); -- sfix8_En12
  CONSTANT coeff278                       : signed(7 DOWNTO 0) := to_signed(-17, 8); -- sfix8_En12
  CONSTANT coeff279                       : signed(7 DOWNTO 0) := to_signed(-17, 8); -- sfix8_En12
  CONSTANT coeff280                       : signed(7 DOWNTO 0) := to_signed(-17, 8); -- sfix8_En12
  CONSTANT coeff281                       : signed(7 DOWNTO 0) := to_signed(-17, 8); -- sfix8_En12
  CONSTANT coeff282                       : signed(7 DOWNTO 0) := to_signed(-17, 8); -- sfix8_En12
  CONSTANT coeff283                       : signed(7 DOWNTO 0) := to_signed(-17, 8); -- sfix8_En12
  CONSTANT coeff284                       : signed(7 DOWNTO 0) := to_signed(-16, 8); -- sfix8_En12
  CONSTANT coeff285                       : signed(7 DOWNTO 0) := to_signed(-16, 8); -- sfix8_En12
  CONSTANT coeff286                       : signed(7 DOWNTO 0) := to_signed(-15, 8); -- sfix8_En12
  CONSTANT coeff287                       : signed(7 DOWNTO 0) := to_signed(-14, 8); -- sfix8_En12
  CONSTANT coeff288                       : signed(7 DOWNTO 0) := to_signed(-14, 8); -- sfix8_En12
  CONSTANT coeff289                       : signed(7 DOWNTO 0) := to_signed(-13, 8); -- sfix8_En12
  CONSTANT coeff290                       : signed(7 DOWNTO 0) := to_signed(-12, 8); -- sfix8_En12
  CONSTANT coeff291                       : signed(7 DOWNTO 0) := to_signed(-11, 8); -- sfix8_En12
  CONSTANT coeff292                       : signed(7 DOWNTO 0) := to_signed(-10, 8); -- sfix8_En12
  CONSTANT coeff293                       : signed(7 DOWNTO 0) := to_signed(-9, 8); -- sfix8_En12
  CONSTANT coeff294                       : signed(7 DOWNTO 0) := to_signed(-8, 8); -- sfix8_En12
  CONSTANT coeff295                       : signed(7 DOWNTO 0) := to_signed(-6, 8); -- sfix8_En12
  CONSTANT coeff296                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff297                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff298                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff299                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff300                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff301                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff302                       : signed(7 DOWNTO 0) := to_signed(5, 8); -- sfix8_En12
  CONSTANT coeff303                       : signed(7 DOWNTO 0) := to_signed(7, 8); -- sfix8_En12
  CONSTANT coeff304                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff305                       : signed(7 DOWNTO 0) := to_signed(11, 8); -- sfix8_En12
  CONSTANT coeff306                       : signed(7 DOWNTO 0) := to_signed(13, 8); -- sfix8_En12
  CONSTANT coeff307                       : signed(7 DOWNTO 0) := to_signed(15, 8); -- sfix8_En12
  CONSTANT coeff308                       : signed(7 DOWNTO 0) := to_signed(18, 8); -- sfix8_En12
  CONSTANT coeff309                       : signed(7 DOWNTO 0) := to_signed(20, 8); -- sfix8_En12
  CONSTANT coeff310                       : signed(7 DOWNTO 0) := to_signed(22, 8); -- sfix8_En12
  CONSTANT coeff311                       : signed(7 DOWNTO 0) := to_signed(24, 8); -- sfix8_En12
  CONSTANT coeff312                       : signed(7 DOWNTO 0) := to_signed(27, 8); -- sfix8_En12
  CONSTANT coeff313                       : signed(7 DOWNTO 0) := to_signed(29, 8); -- sfix8_En12
  CONSTANT coeff314                       : signed(7 DOWNTO 0) := to_signed(32, 8); -- sfix8_En12
  CONSTANT coeff315                       : signed(7 DOWNTO 0) := to_signed(34, 8); -- sfix8_En12
  CONSTANT coeff316                       : signed(7 DOWNTO 0) := to_signed(36, 8); -- sfix8_En12
  CONSTANT coeff317                       : signed(7 DOWNTO 0) := to_signed(39, 8); -- sfix8_En12
  CONSTANT coeff318                       : signed(7 DOWNTO 0) := to_signed(41, 8); -- sfix8_En12
  CONSTANT coeff319                       : signed(7 DOWNTO 0) := to_signed(43, 8); -- sfix8_En12
  CONSTANT coeff320                       : signed(7 DOWNTO 0) := to_signed(46, 8); -- sfix8_En12
  CONSTANT coeff321                       : signed(7 DOWNTO 0) := to_signed(48, 8); -- sfix8_En12
  CONSTANT coeff322                       : signed(7 DOWNTO 0) := to_signed(50, 8); -- sfix8_En12
  CONSTANT coeff323                       : signed(7 DOWNTO 0) := to_signed(53, 8); -- sfix8_En12
  CONSTANT coeff324                       : signed(7 DOWNTO 0) := to_signed(55, 8); -- sfix8_En12
  CONSTANT coeff325                       : signed(7 DOWNTO 0) := to_signed(57, 8); -- sfix8_En12
  CONSTANT coeff326                       : signed(7 DOWNTO 0) := to_signed(59, 8); -- sfix8_En12
  CONSTANT coeff327                       : signed(7 DOWNTO 0) := to_signed(61, 8); -- sfix8_En12
  CONSTANT coeff328                       : signed(7 DOWNTO 0) := to_signed(63, 8); -- sfix8_En12
  CONSTANT coeff329                       : signed(7 DOWNTO 0) := to_signed(65, 8); -- sfix8_En12
  CONSTANT coeff330                       : signed(7 DOWNTO 0) := to_signed(67, 8); -- sfix8_En12
  CONSTANT coeff331                       : signed(7 DOWNTO 0) := to_signed(69, 8); -- sfix8_En12
  CONSTANT coeff332                       : signed(7 DOWNTO 0) := to_signed(71, 8); -- sfix8_En12
  CONSTANT coeff333                       : signed(7 DOWNTO 0) := to_signed(72, 8); -- sfix8_En12
  CONSTANT coeff334                       : signed(7 DOWNTO 0) := to_signed(74, 8); -- sfix8_En12
  CONSTANT coeff335                       : signed(7 DOWNTO 0) := to_signed(75, 8); -- sfix8_En12
  CONSTANT coeff336                       : signed(7 DOWNTO 0) := to_signed(77, 8); -- sfix8_En12
  CONSTANT coeff337                       : signed(7 DOWNTO 0) := to_signed(78, 8); -- sfix8_En12
  CONSTANT coeff338                       : signed(7 DOWNTO 0) := to_signed(79, 8); -- sfix8_En12
  CONSTANT coeff339                       : signed(7 DOWNTO 0) := to_signed(80, 8); -- sfix8_En12
  CONSTANT coeff340                       : signed(7 DOWNTO 0) := to_signed(81, 8); -- sfix8_En12
  CONSTANT coeff341                       : signed(7 DOWNTO 0) := to_signed(82, 8); -- sfix8_En12
  CONSTANT coeff342                       : signed(7 DOWNTO 0) := to_signed(83, 8); -- sfix8_En12
  CONSTANT coeff343                       : signed(7 DOWNTO 0) := to_signed(83, 8); -- sfix8_En12
  CONSTANT coeff344                       : signed(7 DOWNTO 0) := to_signed(84, 8); -- sfix8_En12
  CONSTANT coeff345                       : signed(7 DOWNTO 0) := to_signed(84, 8); -- sfix8_En12
  CONSTANT coeff346                       : signed(7 DOWNTO 0) := to_signed(84, 8); -- sfix8_En12
  CONSTANT coeff347                       : signed(7 DOWNTO 0) := to_signed(85, 8); -- sfix8_En12
  CONSTANT coeff348                       : signed(7 DOWNTO 0) := to_signed(85, 8); -- sfix8_En12
  CONSTANT coeff349                       : signed(7 DOWNTO 0) := to_signed(84, 8); -- sfix8_En12
  CONSTANT coeff350                       : signed(7 DOWNTO 0) := to_signed(84, 8); -- sfix8_En12
  CONSTANT coeff351                       : signed(7 DOWNTO 0) := to_signed(84, 8); -- sfix8_En12
  CONSTANT coeff352                       : signed(7 DOWNTO 0) := to_signed(83, 8); -- sfix8_En12
  CONSTANT coeff353                       : signed(7 DOWNTO 0) := to_signed(83, 8); -- sfix8_En12
  CONSTANT coeff354                       : signed(7 DOWNTO 0) := to_signed(82, 8); -- sfix8_En12
  CONSTANT coeff355                       : signed(7 DOWNTO 0) := to_signed(81, 8); -- sfix8_En12
  CONSTANT coeff356                       : signed(7 DOWNTO 0) := to_signed(80, 8); -- sfix8_En12
  CONSTANT coeff357                       : signed(7 DOWNTO 0) := to_signed(79, 8); -- sfix8_En12
  CONSTANT coeff358                       : signed(7 DOWNTO 0) := to_signed(78, 8); -- sfix8_En12
  CONSTANT coeff359                       : signed(7 DOWNTO 0) := to_signed(77, 8); -- sfix8_En12
  CONSTANT coeff360                       : signed(7 DOWNTO 0) := to_signed(75, 8); -- sfix8_En12
  CONSTANT coeff361                       : signed(7 DOWNTO 0) := to_signed(74, 8); -- sfix8_En12
  CONSTANT coeff362                       : signed(7 DOWNTO 0) := to_signed(72, 8); -- sfix8_En12
  CONSTANT coeff363                       : signed(7 DOWNTO 0) := to_signed(71, 8); -- sfix8_En12
  CONSTANT coeff364                       : signed(7 DOWNTO 0) := to_signed(69, 8); -- sfix8_En12
  CONSTANT coeff365                       : signed(7 DOWNTO 0) := to_signed(67, 8); -- sfix8_En12
  CONSTANT coeff366                       : signed(7 DOWNTO 0) := to_signed(65, 8); -- sfix8_En12
  CONSTANT coeff367                       : signed(7 DOWNTO 0) := to_signed(63, 8); -- sfix8_En12
  CONSTANT coeff368                       : signed(7 DOWNTO 0) := to_signed(61, 8); -- sfix8_En12
  CONSTANT coeff369                       : signed(7 DOWNTO 0) := to_signed(59, 8); -- sfix8_En12
  CONSTANT coeff370                       : signed(7 DOWNTO 0) := to_signed(57, 8); -- sfix8_En12
  CONSTANT coeff371                       : signed(7 DOWNTO 0) := to_signed(55, 8); -- sfix8_En12
  CONSTANT coeff372                       : signed(7 DOWNTO 0) := to_signed(53, 8); -- sfix8_En12
  CONSTANT coeff373                       : signed(7 DOWNTO 0) := to_signed(50, 8); -- sfix8_En12
  CONSTANT coeff374                       : signed(7 DOWNTO 0) := to_signed(48, 8); -- sfix8_En12
  CONSTANT coeff375                       : signed(7 DOWNTO 0) := to_signed(46, 8); -- sfix8_En12
  CONSTANT coeff376                       : signed(7 DOWNTO 0) := to_signed(43, 8); -- sfix8_En12
  CONSTANT coeff377                       : signed(7 DOWNTO 0) := to_signed(41, 8); -- sfix8_En12
  CONSTANT coeff378                       : signed(7 DOWNTO 0) := to_signed(39, 8); -- sfix8_En12
  CONSTANT coeff379                       : signed(7 DOWNTO 0) := to_signed(36, 8); -- sfix8_En12
  CONSTANT coeff380                       : signed(7 DOWNTO 0) := to_signed(34, 8); -- sfix8_En12
  CONSTANT coeff381                       : signed(7 DOWNTO 0) := to_signed(32, 8); -- sfix8_En12
  CONSTANT coeff382                       : signed(7 DOWNTO 0) := to_signed(29, 8); -- sfix8_En12
  CONSTANT coeff383                       : signed(7 DOWNTO 0) := to_signed(27, 8); -- sfix8_En12
  CONSTANT coeff384                       : signed(7 DOWNTO 0) := to_signed(24, 8); -- sfix8_En12
  CONSTANT coeff385                       : signed(7 DOWNTO 0) := to_signed(22, 8); -- sfix8_En12
  CONSTANT coeff386                       : signed(7 DOWNTO 0) := to_signed(20, 8); -- sfix8_En12
  CONSTANT coeff387                       : signed(7 DOWNTO 0) := to_signed(18, 8); -- sfix8_En12
  CONSTANT coeff388                       : signed(7 DOWNTO 0) := to_signed(15, 8); -- sfix8_En12
  CONSTANT coeff389                       : signed(7 DOWNTO 0) := to_signed(13, 8); -- sfix8_En12
  CONSTANT coeff390                       : signed(7 DOWNTO 0) := to_signed(11, 8); -- sfix8_En12
  CONSTANT coeff391                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff392                       : signed(7 DOWNTO 0) := to_signed(7, 8); -- sfix8_En12
  CONSTANT coeff393                       : signed(7 DOWNTO 0) := to_signed(5, 8); -- sfix8_En12
  CONSTANT coeff394                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff395                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff396                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff397                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff398                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff399                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff400                       : signed(7 DOWNTO 0) := to_signed(-6, 8); -- sfix8_En12
  CONSTANT coeff401                       : signed(7 DOWNTO 0) := to_signed(-8, 8); -- sfix8_En12
  CONSTANT coeff402                       : signed(7 DOWNTO 0) := to_signed(-9, 8); -- sfix8_En12
  CONSTANT coeff403                       : signed(7 DOWNTO 0) := to_signed(-10, 8); -- sfix8_En12
  CONSTANT coeff404                       : signed(7 DOWNTO 0) := to_signed(-11, 8); -- sfix8_En12
  CONSTANT coeff405                       : signed(7 DOWNTO 0) := to_signed(-12, 8); -- sfix8_En12
  CONSTANT coeff406                       : signed(7 DOWNTO 0) := to_signed(-13, 8); -- sfix8_En12
  CONSTANT coeff407                       : signed(7 DOWNTO 0) := to_signed(-14, 8); -- sfix8_En12
  CONSTANT coeff408                       : signed(7 DOWNTO 0) := to_signed(-14, 8); -- sfix8_En12
  CONSTANT coeff409                       : signed(7 DOWNTO 0) := to_signed(-15, 8); -- sfix8_En12
  CONSTANT coeff410                       : signed(7 DOWNTO 0) := to_signed(-16, 8); -- sfix8_En12
  CONSTANT coeff411                       : signed(7 DOWNTO 0) := to_signed(-16, 8); -- sfix8_En12
  CONSTANT coeff412                       : signed(7 DOWNTO 0) := to_signed(-17, 8); -- sfix8_En12
  CONSTANT coeff413                       : signed(7 DOWNTO 0) := to_signed(-17, 8); -- sfix8_En12
  CONSTANT coeff414                       : signed(7 DOWNTO 0) := to_signed(-17, 8); -- sfix8_En12
  CONSTANT coeff415                       : signed(7 DOWNTO 0) := to_signed(-17, 8); -- sfix8_En12
  CONSTANT coeff416                       : signed(7 DOWNTO 0) := to_signed(-17, 8); -- sfix8_En12
  CONSTANT coeff417                       : signed(7 DOWNTO 0) := to_signed(-17, 8); -- sfix8_En12
  CONSTANT coeff418                       : signed(7 DOWNTO 0) := to_signed(-17, 8); -- sfix8_En12
  CONSTANT coeff419                       : signed(7 DOWNTO 0) := to_signed(-17, 8); -- sfix8_En12
  CONSTANT coeff420                       : signed(7 DOWNTO 0) := to_signed(-17, 8); -- sfix8_En12
  CONSTANT coeff421                       : signed(7 DOWNTO 0) := to_signed(-16, 8); -- sfix8_En12
  CONSTANT coeff422                       : signed(7 DOWNTO 0) := to_signed(-16, 8); -- sfix8_En12
  CONSTANT coeff423                       : signed(7 DOWNTO 0) := to_signed(-16, 8); -- sfix8_En12
  CONSTANT coeff424                       : signed(7 DOWNTO 0) := to_signed(-15, 8); -- sfix8_En12
  CONSTANT coeff425                       : signed(7 DOWNTO 0) := to_signed(-15, 8); -- sfix8_En12
  CONSTANT coeff426                       : signed(7 DOWNTO 0) := to_signed(-14, 8); -- sfix8_En12
  CONSTANT coeff427                       : signed(7 DOWNTO 0) := to_signed(-14, 8); -- sfix8_En12
  CONSTANT coeff428                       : signed(7 DOWNTO 0) := to_signed(-13, 8); -- sfix8_En12
  CONSTANT coeff429                       : signed(7 DOWNTO 0) := to_signed(-12, 8); -- sfix8_En12
  CONSTANT coeff430                       : signed(7 DOWNTO 0) := to_signed(-11, 8); -- sfix8_En12
  CONSTANT coeff431                       : signed(7 DOWNTO 0) := to_signed(-11, 8); -- sfix8_En12
  CONSTANT coeff432                       : signed(7 DOWNTO 0) := to_signed(-10, 8); -- sfix8_En12
  CONSTANT coeff433                       : signed(7 DOWNTO 0) := to_signed(-9, 8); -- sfix8_En12
  CONSTANT coeff434                       : signed(7 DOWNTO 0) := to_signed(-8, 8); -- sfix8_En12
  CONSTANT coeff435                       : signed(7 DOWNTO 0) := to_signed(-8, 8); -- sfix8_En12
  CONSTANT coeff436                       : signed(7 DOWNTO 0) := to_signed(-7, 8); -- sfix8_En12
  CONSTANT coeff437                       : signed(7 DOWNTO 0) := to_signed(-6, 8); -- sfix8_En12
  CONSTANT coeff438                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff439                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff440                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff441                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff442                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff443                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff444                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff445                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff446                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff447                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff448                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff449                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff450                       : signed(7 DOWNTO 0) := to_signed(4, 8); -- sfix8_En12
  CONSTANT coeff451                       : signed(7 DOWNTO 0) := to_signed(5, 8); -- sfix8_En12
  CONSTANT coeff452                       : signed(7 DOWNTO 0) := to_signed(5, 8); -- sfix8_En12
  CONSTANT coeff453                       : signed(7 DOWNTO 0) := to_signed(6, 8); -- sfix8_En12
  CONSTANT coeff454                       : signed(7 DOWNTO 0) := to_signed(6, 8); -- sfix8_En12
  CONSTANT coeff455                       : signed(7 DOWNTO 0) := to_signed(7, 8); -- sfix8_En12
  CONSTANT coeff456                       : signed(7 DOWNTO 0) := to_signed(7, 8); -- sfix8_En12
  CONSTANT coeff457                       : signed(7 DOWNTO 0) := to_signed(7, 8); -- sfix8_En12
  CONSTANT coeff458                       : signed(7 DOWNTO 0) := to_signed(8, 8); -- sfix8_En12
  CONSTANT coeff459                       : signed(7 DOWNTO 0) := to_signed(8, 8); -- sfix8_En12
  CONSTANT coeff460                       : signed(7 DOWNTO 0) := to_signed(8, 8); -- sfix8_En12
  CONSTANT coeff461                       : signed(7 DOWNTO 0) := to_signed(8, 8); -- sfix8_En12
  CONSTANT coeff462                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff463                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff464                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff465                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff466                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff467                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff468                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff469                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff470                       : signed(7 DOWNTO 0) := to_signed(9, 8); -- sfix8_En12
  CONSTANT coeff471                       : signed(7 DOWNTO 0) := to_signed(8, 8); -- sfix8_En12
  CONSTANT coeff472                       : signed(7 DOWNTO 0) := to_signed(8, 8); -- sfix8_En12
  CONSTANT coeff473                       : signed(7 DOWNTO 0) := to_signed(8, 8); -- sfix8_En12
  CONSTANT coeff474                       : signed(7 DOWNTO 0) := to_signed(8, 8); -- sfix8_En12
  CONSTANT coeff475                       : signed(7 DOWNTO 0) := to_signed(7, 8); -- sfix8_En12
  CONSTANT coeff476                       : signed(7 DOWNTO 0) := to_signed(7, 8); -- sfix8_En12
  CONSTANT coeff477                       : signed(7 DOWNTO 0) := to_signed(7, 8); -- sfix8_En12
  CONSTANT coeff478                       : signed(7 DOWNTO 0) := to_signed(6, 8); -- sfix8_En12
  CONSTANT coeff479                       : signed(7 DOWNTO 0) := to_signed(6, 8); -- sfix8_En12
  CONSTANT coeff480                       : signed(7 DOWNTO 0) := to_signed(6, 8); -- sfix8_En12
  CONSTANT coeff481                       : signed(7 DOWNTO 0) := to_signed(5, 8); -- sfix8_En12
  CONSTANT coeff482                       : signed(7 DOWNTO 0) := to_signed(5, 8); -- sfix8_En12
  CONSTANT coeff483                       : signed(7 DOWNTO 0) := to_signed(4, 8); -- sfix8_En12
  CONSTANT coeff484                       : signed(7 DOWNTO 0) := to_signed(4, 8); -- sfix8_En12
  CONSTANT coeff485                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff486                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff487                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff488                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff489                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff490                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff491                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff492                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff493                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff494                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff495                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff496                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff497                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff498                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff499                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff500                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff501                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff502                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff503                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff504                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff505                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff506                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff507                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff508                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff509                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff510                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff511                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff512                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff513                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff514                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff515                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff516                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff517                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff518                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff519                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff520                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff521                       : signed(7 DOWNTO 0) := to_signed(-5, 8); -- sfix8_En12
  CONSTANT coeff522                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff523                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff524                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff525                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff526                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff527                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff528                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff529                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff530                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff531                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff532                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff533                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff534                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff535                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff536                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff537                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff538                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff539                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff540                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff541                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff542                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff543                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff544                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff545                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff546                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff547                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff548                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff549                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff550                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff551                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff552                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff553                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff554                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff555                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff556                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff557                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff558                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff559                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff560                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff561                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff562                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff563                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff564                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff565                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff566                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff567                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff568                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff569                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff570                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff571                       : signed(7 DOWNTO 0) := to_signed(3, 8); -- sfix8_En12
  CONSTANT coeff572                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff573                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff574                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff575                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff576                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff577                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff578                       : signed(7 DOWNTO 0) := to_signed(2, 8); -- sfix8_En12
  CONSTANT coeff579                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff580                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff581                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff582                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff583                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff584                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff585                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff586                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff587                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff588                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff589                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff590                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff591                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff592                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff593                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff594                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff595                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff596                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff597                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff598                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff599                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff600                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff601                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff602                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff603                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff604                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff605                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff606                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff607                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff608                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff609                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff610                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff611                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff612                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff613                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff614                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff615                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff616                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff617                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff618                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff619                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff620                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff621                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff622                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff623                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff624                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff625                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff626                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff627                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff628                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff629                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff630                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff631                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff632                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff633                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff634                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff635                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff636                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff637                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff638                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff639                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff640                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff641                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff642                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff643                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff644                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff645                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff646                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff647                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff648                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff649                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff650                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff651                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff652                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff653                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff654                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff655                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff656                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff657                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff658                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff659                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff660                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff661                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff662                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff663                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff664                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff665                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff666                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff667                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff668                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff669                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff670                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff671                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff672                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff673                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff674                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff675                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff676                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff677                       : signed(7 DOWNTO 0) := to_signed(1, 8); -- sfix8_En12
  CONSTANT coeff678                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff679                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff680                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff681                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff682                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff683                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff684                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff685                       : signed(7 DOWNTO 0) := to_signed(0, 8); -- sfix8_En12
  CONSTANT coeff686                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff687                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff688                       : signed(7 DOWNTO 0) := to_signed(-1, 8); -- sfix8_En12
  CONSTANT coeff689                       : signed(7 DOWNTO 0) := to_signed(-2, 8); -- sfix8_En12
  CONSTANT coeff690                       : signed(7 DOWNTO 0) := to_signed(-3, 8); -- sfix8_En12
  CONSTANT coeff691                       : signed(7 DOWNTO 0) := to_signed(-4, 8); -- sfix8_En12
  CONSTANT coeff692                       : signed(7 DOWNTO 0) := to_signed(-6, 8); -- sfix8_En12
  CONSTANT coeff693                       : signed(7 DOWNTO 0) := to_signed(-8, 8); -- sfix8_En12
  CONSTANT coeff694                       : signed(7 DOWNTO 0) := to_signed(13, 8); -- sfix8_En12

  -- Signals
  SIGNAL cur_count                        : unsigned(9 DOWNTO 0); -- ufix10
  SIGNAL phase_0                          : std_logic; -- boolean
  SIGNAL delay_pipeline                   : delay_pipeline_type(0 TO 693); -- sfix32_En31
  SIGNAL I_FILTER_regtype                 : signed(31 DOWNTO 0); -- sfix32_En31
  SIGNAL inputmux_1                       : signed(31 DOWNTO 0); -- sfix32_En31
  SIGNAL acc_final                        : signed(44 DOWNTO 0); -- sfix45_En43
  SIGNAL acc_out_1                        : signed(44 DOWNTO 0); -- sfix45_En43
  SIGNAL product_1                        : signed(38 DOWNTO 0); -- sfix39_En43
  SIGNAL product_1_mux                    : signed(7 DOWNTO 0); -- sfix8_En12
  SIGNAL mul_temp                         : signed(39 DOWNTO 0); -- sfix40_En43
  SIGNAL prod_typeconvert_1               : signed(44 DOWNTO 0); -- sfix45_En43
  SIGNAL acc_sum_1                        : signed(44 DOWNTO 0); -- sfix45_En43
  SIGNAL acc_in_1                         : signed(44 DOWNTO 0); -- sfix45_En43
  SIGNAL add_temp                         : signed(45 DOWNTO 0); -- sfix46_En43
  SIGNAL output_typeconvert               : signed(44 DOWNTO 0); -- sfix45_En43
  SIGNAL output_register                  : signed(44 DOWNTO 0); -- sfix45_En43


BEGIN

  -- Block Statements
  Counter_process : PROCESS (I_CLK, I_RST)
  BEGIN
    IF I_RST = '1' THEN
      cur_count <= to_unsigned(0, 10);
    ELSIF rising_edge(I_CLK) THEN
      IF cur_count >= to_unsigned(621, 10) THEN
        cur_count <= to_unsigned(0, 10);
      ELSE
        cur_count <= cur_count + to_unsigned(1, 10);
      END IF;
    END IF;
  END PROCESS Counter_process;

  phase_0 <= '1' WHEN cur_count = to_unsigned(0, 10) ELSE '0';

  Delay_Pipeline_process : PROCESS (I_CLK, I_RST)
  BEGIN
    IF I_RST = '1' THEN
      delay_pipeline(0 TO 693) <= (OTHERS => (OTHERS => '0'));
    ELSIF rising_edge(I_CLK) THEN
      IF phase_0 = '1' THEN
        delay_pipeline(0) <= signed(I_FILTER);
        delay_pipeline(1 TO 693) <= delay_pipeline(0 TO 692);
      END IF;
    END IF;
  END PROCESS Delay_Pipeline_process;

  I_FILTER_regtype <= signed(I_FILTER);

  inputmux_1 <= I_FILTER_regtype WHEN ( cur_count = to_unsigned(0, 10) ) ELSE
                     delay_pipeline(1) WHEN ( cur_count = to_unsigned(1, 10) ) ELSE
                     delay_pipeline(2) WHEN ( cur_count = to_unsigned(2, 10) ) ELSE
                     delay_pipeline(3) WHEN ( cur_count = to_unsigned(3, 10) ) ELSE
                     delay_pipeline(4) WHEN ( cur_count = to_unsigned(4, 10) ) ELSE
                     delay_pipeline(5) WHEN ( cur_count = to_unsigned(5, 10) ) ELSE
                     delay_pipeline(6) WHEN ( cur_count = to_unsigned(6, 10) ) ELSE
                     delay_pipeline(7) WHEN ( cur_count = to_unsigned(7, 10) ) ELSE
                     delay_pipeline(8) WHEN ( cur_count = to_unsigned(8, 10) ) ELSE
                     delay_pipeline(17) WHEN ( cur_count = to_unsigned(9, 10) ) ELSE
                     delay_pipeline(18) WHEN ( cur_count = to_unsigned(10, 10) ) ELSE
                     delay_pipeline(19) WHEN ( cur_count = to_unsigned(11, 10) ) ELSE
                     delay_pipeline(20) WHEN ( cur_count = to_unsigned(12, 10) ) ELSE
                     delay_pipeline(21) WHEN ( cur_count = to_unsigned(13, 10) ) ELSE
                     delay_pipeline(22) WHEN ( cur_count = to_unsigned(14, 10) ) ELSE
                     delay_pipeline(23) WHEN ( cur_count = to_unsigned(15, 10) ) ELSE
                     delay_pipeline(24) WHEN ( cur_count = to_unsigned(16, 10) ) ELSE
                     delay_pipeline(25) WHEN ( cur_count = to_unsigned(17, 10) ) ELSE
                     delay_pipeline(26) WHEN ( cur_count = to_unsigned(18, 10) ) ELSE
                     delay_pipeline(27) WHEN ( cur_count = to_unsigned(19, 10) ) ELSE
                     delay_pipeline(28) WHEN ( cur_count = to_unsigned(20, 10) ) ELSE
                     delay_pipeline(29) WHEN ( cur_count = to_unsigned(21, 10) ) ELSE
                     delay_pipeline(30) WHEN ( cur_count = to_unsigned(22, 10) ) ELSE
                     delay_pipeline(31) WHEN ( cur_count = to_unsigned(23, 10) ) ELSE
                     delay_pipeline(32) WHEN ( cur_count = to_unsigned(24, 10) ) ELSE
                     delay_pipeline(33) WHEN ( cur_count = to_unsigned(25, 10) ) ELSE
                     delay_pipeline(34) WHEN ( cur_count = to_unsigned(26, 10) ) ELSE
                     delay_pipeline(35) WHEN ( cur_count = to_unsigned(27, 10) ) ELSE
                     delay_pipeline(36) WHEN ( cur_count = to_unsigned(28, 10) ) ELSE
                     delay_pipeline(37) WHEN ( cur_count = to_unsigned(29, 10) ) ELSE
                     delay_pipeline(38) WHEN ( cur_count = to_unsigned(30, 10) ) ELSE
                     delay_pipeline(39) WHEN ( cur_count = to_unsigned(31, 10) ) ELSE
                     delay_pipeline(40) WHEN ( cur_count = to_unsigned(32, 10) ) ELSE
                     delay_pipeline(41) WHEN ( cur_count = to_unsigned(33, 10) ) ELSE
                     delay_pipeline(42) WHEN ( cur_count = to_unsigned(34, 10) ) ELSE
                     delay_pipeline(43) WHEN ( cur_count = to_unsigned(35, 10) ) ELSE
                     delay_pipeline(44) WHEN ( cur_count = to_unsigned(36, 10) ) ELSE
                     delay_pipeline(45) WHEN ( cur_count = to_unsigned(37, 10) ) ELSE
                     delay_pipeline(46) WHEN ( cur_count = to_unsigned(38, 10) ) ELSE
                     delay_pipeline(47) WHEN ( cur_count = to_unsigned(39, 10) ) ELSE
                     delay_pipeline(48) WHEN ( cur_count = to_unsigned(40, 10) ) ELSE
                     delay_pipeline(49) WHEN ( cur_count = to_unsigned(41, 10) ) ELSE
                     delay_pipeline(50) WHEN ( cur_count = to_unsigned(42, 10) ) ELSE
                     delay_pipeline(51) WHEN ( cur_count = to_unsigned(43, 10) ) ELSE
                     delay_pipeline(65) WHEN ( cur_count = to_unsigned(44, 10) ) ELSE
                     delay_pipeline(66) WHEN ( cur_count = to_unsigned(45, 10) ) ELSE
                     delay_pipeline(67) WHEN ( cur_count = to_unsigned(46, 10) ) ELSE
                     delay_pipeline(68) WHEN ( cur_count = to_unsigned(47, 10) ) ELSE
                     delay_pipeline(69) WHEN ( cur_count = to_unsigned(48, 10) ) ELSE
                     delay_pipeline(70) WHEN ( cur_count = to_unsigned(49, 10) ) ELSE
                     delay_pipeline(71) WHEN ( cur_count = to_unsigned(50, 10) ) ELSE
                     delay_pipeline(72) WHEN ( cur_count = to_unsigned(51, 10) ) ELSE
                     delay_pipeline(73) WHEN ( cur_count = to_unsigned(52, 10) ) ELSE
                     delay_pipeline(74) WHEN ( cur_count = to_unsigned(53, 10) ) ELSE
                     delay_pipeline(75) WHEN ( cur_count = to_unsigned(54, 10) ) ELSE
                     delay_pipeline(76) WHEN ( cur_count = to_unsigned(55, 10) ) ELSE
                     delay_pipeline(77) WHEN ( cur_count = to_unsigned(56, 10) ) ELSE
                     delay_pipeline(78) WHEN ( cur_count = to_unsigned(57, 10) ) ELSE
                     delay_pipeline(79) WHEN ( cur_count = to_unsigned(58, 10) ) ELSE
                     delay_pipeline(80) WHEN ( cur_count = to_unsigned(59, 10) ) ELSE
                     delay_pipeline(81) WHEN ( cur_count = to_unsigned(60, 10) ) ELSE
                     delay_pipeline(82) WHEN ( cur_count = to_unsigned(61, 10) ) ELSE
                     delay_pipeline(83) WHEN ( cur_count = to_unsigned(62, 10) ) ELSE
                     delay_pipeline(84) WHEN ( cur_count = to_unsigned(63, 10) ) ELSE
                     delay_pipeline(85) WHEN ( cur_count = to_unsigned(64, 10) ) ELSE
                     delay_pipeline(86) WHEN ( cur_count = to_unsigned(65, 10) ) ELSE
                     delay_pipeline(87) WHEN ( cur_count = to_unsigned(66, 10) ) ELSE
                     delay_pipeline(88) WHEN ( cur_count = to_unsigned(67, 10) ) ELSE
                     delay_pipeline(89) WHEN ( cur_count = to_unsigned(68, 10) ) ELSE
                     delay_pipeline(90) WHEN ( cur_count = to_unsigned(69, 10) ) ELSE
                     delay_pipeline(91) WHEN ( cur_count = to_unsigned(70, 10) ) ELSE
                     delay_pipeline(92) WHEN ( cur_count = to_unsigned(71, 10) ) ELSE
                     delay_pipeline(93) WHEN ( cur_count = to_unsigned(72, 10) ) ELSE
                     delay_pipeline(94) WHEN ( cur_count = to_unsigned(73, 10) ) ELSE
                     delay_pipeline(95) WHEN ( cur_count = to_unsigned(74, 10) ) ELSE
                     delay_pipeline(96) WHEN ( cur_count = to_unsigned(75, 10) ) ELSE
                     delay_pipeline(97) WHEN ( cur_count = to_unsigned(76, 10) ) ELSE
                     delay_pipeline(98) WHEN ( cur_count = to_unsigned(77, 10) ) ELSE
                     delay_pipeline(99) WHEN ( cur_count = to_unsigned(78, 10) ) ELSE
                     delay_pipeline(100) WHEN ( cur_count = to_unsigned(79, 10) ) ELSE
                     delay_pipeline(101) WHEN ( cur_count = to_unsigned(80, 10) ) ELSE
                     delay_pipeline(102) WHEN ( cur_count = to_unsigned(81, 10) ) ELSE
                     delay_pipeline(110) WHEN ( cur_count = to_unsigned(82, 10) ) ELSE
                     delay_pipeline(111) WHEN ( cur_count = to_unsigned(83, 10) ) ELSE
                     delay_pipeline(112) WHEN ( cur_count = to_unsigned(84, 10) ) ELSE
                     delay_pipeline(113) WHEN ( cur_count = to_unsigned(85, 10) ) ELSE
                     delay_pipeline(114) WHEN ( cur_count = to_unsigned(86, 10) ) ELSE
                     delay_pipeline(115) WHEN ( cur_count = to_unsigned(87, 10) ) ELSE
                     delay_pipeline(116) WHEN ( cur_count = to_unsigned(88, 10) ) ELSE
                     delay_pipeline(117) WHEN ( cur_count = to_unsigned(89, 10) ) ELSE
                     delay_pipeline(118) WHEN ( cur_count = to_unsigned(90, 10) ) ELSE
                     delay_pipeline(119) WHEN ( cur_count = to_unsigned(91, 10) ) ELSE
                     delay_pipeline(120) WHEN ( cur_count = to_unsigned(92, 10) ) ELSE
                     delay_pipeline(121) WHEN ( cur_count = to_unsigned(93, 10) ) ELSE
                     delay_pipeline(122) WHEN ( cur_count = to_unsigned(94, 10) ) ELSE
                     delay_pipeline(123) WHEN ( cur_count = to_unsigned(95, 10) ) ELSE
                     delay_pipeline(124) WHEN ( cur_count = to_unsigned(96, 10) ) ELSE
                     delay_pipeline(125) WHEN ( cur_count = to_unsigned(97, 10) ) ELSE
                     delay_pipeline(126) WHEN ( cur_count = to_unsigned(98, 10) ) ELSE
                     delay_pipeline(127) WHEN ( cur_count = to_unsigned(99, 10) ) ELSE
                     delay_pipeline(128) WHEN ( cur_count = to_unsigned(100, 10) ) ELSE
                     delay_pipeline(129) WHEN ( cur_count = to_unsigned(101, 10) ) ELSE
                     delay_pipeline(130) WHEN ( cur_count = to_unsigned(102, 10) ) ELSE
                     delay_pipeline(131) WHEN ( cur_count = to_unsigned(103, 10) ) ELSE
                     delay_pipeline(132) WHEN ( cur_count = to_unsigned(104, 10) ) ELSE
                     delay_pipeline(133) WHEN ( cur_count = to_unsigned(105, 10) ) ELSE
                     delay_pipeline(134) WHEN ( cur_count = to_unsigned(106, 10) ) ELSE
                     delay_pipeline(135) WHEN ( cur_count = to_unsigned(107, 10) ) ELSE
                     delay_pipeline(136) WHEN ( cur_count = to_unsigned(108, 10) ) ELSE
                     delay_pipeline(137) WHEN ( cur_count = to_unsigned(109, 10) ) ELSE
                     delay_pipeline(138) WHEN ( cur_count = to_unsigned(110, 10) ) ELSE
                     delay_pipeline(139) WHEN ( cur_count = to_unsigned(111, 10) ) ELSE
                     delay_pipeline(140) WHEN ( cur_count = to_unsigned(112, 10) ) ELSE
                     delay_pipeline(141) WHEN ( cur_count = to_unsigned(113, 10) ) ELSE
                     delay_pipeline(142) WHEN ( cur_count = to_unsigned(114, 10) ) ELSE
                     delay_pipeline(143) WHEN ( cur_count = to_unsigned(115, 10) ) ELSE
                     delay_pipeline(144) WHEN ( cur_count = to_unsigned(116, 10) ) ELSE
                     delay_pipeline(145) WHEN ( cur_count = to_unsigned(117, 10) ) ELSE
                     delay_pipeline(146) WHEN ( cur_count = to_unsigned(118, 10) ) ELSE
                     delay_pipeline(147) WHEN ( cur_count = to_unsigned(119, 10) ) ELSE
                     delay_pipeline(148) WHEN ( cur_count = to_unsigned(120, 10) ) ELSE
                     delay_pipeline(149) WHEN ( cur_count = to_unsigned(121, 10) ) ELSE
                     delay_pipeline(150) WHEN ( cur_count = to_unsigned(122, 10) ) ELSE
                     delay_pipeline(151) WHEN ( cur_count = to_unsigned(123, 10) ) ELSE
                     delay_pipeline(156) WHEN ( cur_count = to_unsigned(124, 10) ) ELSE
                     delay_pipeline(157) WHEN ( cur_count = to_unsigned(125, 10) ) ELSE
                     delay_pipeline(158) WHEN ( cur_count = to_unsigned(126, 10) ) ELSE
                     delay_pipeline(159) WHEN ( cur_count = to_unsigned(127, 10) ) ELSE
                     delay_pipeline(160) WHEN ( cur_count = to_unsigned(128, 10) ) ELSE
                     delay_pipeline(161) WHEN ( cur_count = to_unsigned(129, 10) ) ELSE
                     delay_pipeline(162) WHEN ( cur_count = to_unsigned(130, 10) ) ELSE
                     delay_pipeline(163) WHEN ( cur_count = to_unsigned(131, 10) ) ELSE
                     delay_pipeline(164) WHEN ( cur_count = to_unsigned(132, 10) ) ELSE
                     delay_pipeline(165) WHEN ( cur_count = to_unsigned(133, 10) ) ELSE
                     delay_pipeline(166) WHEN ( cur_count = to_unsigned(134, 10) ) ELSE
                     delay_pipeline(167) WHEN ( cur_count = to_unsigned(135, 10) ) ELSE
                     delay_pipeline(168) WHEN ( cur_count = to_unsigned(136, 10) ) ELSE
                     delay_pipeline(169) WHEN ( cur_count = to_unsigned(137, 10) ) ELSE
                     delay_pipeline(170) WHEN ( cur_count = to_unsigned(138, 10) ) ELSE
                     delay_pipeline(171) WHEN ( cur_count = to_unsigned(139, 10) ) ELSE
                     delay_pipeline(172) WHEN ( cur_count = to_unsigned(140, 10) ) ELSE
                     delay_pipeline(173) WHEN ( cur_count = to_unsigned(141, 10) ) ELSE
                     delay_pipeline(174) WHEN ( cur_count = to_unsigned(142, 10) ) ELSE
                     delay_pipeline(175) WHEN ( cur_count = to_unsigned(143, 10) ) ELSE
                     delay_pipeline(176) WHEN ( cur_count = to_unsigned(144, 10) ) ELSE
                     delay_pipeline(177) WHEN ( cur_count = to_unsigned(145, 10) ) ELSE
                     delay_pipeline(178) WHEN ( cur_count = to_unsigned(146, 10) ) ELSE
                     delay_pipeline(179) WHEN ( cur_count = to_unsigned(147, 10) ) ELSE
                     delay_pipeline(180) WHEN ( cur_count = to_unsigned(148, 10) ) ELSE
                     delay_pipeline(181) WHEN ( cur_count = to_unsigned(149, 10) ) ELSE
                     delay_pipeline(182) WHEN ( cur_count = to_unsigned(150, 10) ) ELSE
                     delay_pipeline(183) WHEN ( cur_count = to_unsigned(151, 10) ) ELSE
                     delay_pipeline(184) WHEN ( cur_count = to_unsigned(152, 10) ) ELSE
                     delay_pipeline(185) WHEN ( cur_count = to_unsigned(153, 10) ) ELSE
                     delay_pipeline(186) WHEN ( cur_count = to_unsigned(154, 10) ) ELSE
                     delay_pipeline(187) WHEN ( cur_count = to_unsigned(155, 10) ) ELSE
                     delay_pipeline(188) WHEN ( cur_count = to_unsigned(156, 10) ) ELSE
                     delay_pipeline(189) WHEN ( cur_count = to_unsigned(157, 10) ) ELSE
                     delay_pipeline(190) WHEN ( cur_count = to_unsigned(158, 10) ) ELSE
                     delay_pipeline(191) WHEN ( cur_count = to_unsigned(159, 10) ) ELSE
                     delay_pipeline(192) WHEN ( cur_count = to_unsigned(160, 10) ) ELSE
                     delay_pipeline(193) WHEN ( cur_count = to_unsigned(161, 10) ) ELSE
                     delay_pipeline(194) WHEN ( cur_count = to_unsigned(162, 10) ) ELSE
                     delay_pipeline(195) WHEN ( cur_count = to_unsigned(163, 10) ) ELSE
                     delay_pipeline(196) WHEN ( cur_count = to_unsigned(164, 10) ) ELSE
                     delay_pipeline(197) WHEN ( cur_count = to_unsigned(165, 10) ) ELSE
                     delay_pipeline(198) WHEN ( cur_count = to_unsigned(166, 10) ) ELSE
                     delay_pipeline(199) WHEN ( cur_count = to_unsigned(167, 10) ) ELSE
                     delay_pipeline(200) WHEN ( cur_count = to_unsigned(168, 10) ) ELSE
                     delay_pipeline(203) WHEN ( cur_count = to_unsigned(169, 10) ) ELSE
                     delay_pipeline(204) WHEN ( cur_count = to_unsigned(170, 10) ) ELSE
                     delay_pipeline(205) WHEN ( cur_count = to_unsigned(171, 10) ) ELSE
                     delay_pipeline(206) WHEN ( cur_count = to_unsigned(172, 10) ) ELSE
                     delay_pipeline(207) WHEN ( cur_count = to_unsigned(173, 10) ) ELSE
                     delay_pipeline(208) WHEN ( cur_count = to_unsigned(174, 10) ) ELSE
                     delay_pipeline(209) WHEN ( cur_count = to_unsigned(175, 10) ) ELSE
                     delay_pipeline(210) WHEN ( cur_count = to_unsigned(176, 10) ) ELSE
                     delay_pipeline(211) WHEN ( cur_count = to_unsigned(177, 10) ) ELSE
                     delay_pipeline(212) WHEN ( cur_count = to_unsigned(178, 10) ) ELSE
                     delay_pipeline(213) WHEN ( cur_count = to_unsigned(179, 10) ) ELSE
                     delay_pipeline(214) WHEN ( cur_count = to_unsigned(180, 10) ) ELSE
                     delay_pipeline(215) WHEN ( cur_count = to_unsigned(181, 10) ) ELSE
                     delay_pipeline(216) WHEN ( cur_count = to_unsigned(182, 10) ) ELSE
                     delay_pipeline(217) WHEN ( cur_count = to_unsigned(183, 10) ) ELSE
                     delay_pipeline(218) WHEN ( cur_count = to_unsigned(184, 10) ) ELSE
                     delay_pipeline(219) WHEN ( cur_count = to_unsigned(185, 10) ) ELSE
                     delay_pipeline(220) WHEN ( cur_count = to_unsigned(186, 10) ) ELSE
                     delay_pipeline(221) WHEN ( cur_count = to_unsigned(187, 10) ) ELSE
                     delay_pipeline(222) WHEN ( cur_count = to_unsigned(188, 10) ) ELSE
                     delay_pipeline(223) WHEN ( cur_count = to_unsigned(189, 10) ) ELSE
                     delay_pipeline(224) WHEN ( cur_count = to_unsigned(190, 10) ) ELSE
                     delay_pipeline(225) WHEN ( cur_count = to_unsigned(191, 10) ) ELSE
                     delay_pipeline(226) WHEN ( cur_count = to_unsigned(192, 10) ) ELSE
                     delay_pipeline(227) WHEN ( cur_count = to_unsigned(193, 10) ) ELSE
                     delay_pipeline(228) WHEN ( cur_count = to_unsigned(194, 10) ) ELSE
                     delay_pipeline(229) WHEN ( cur_count = to_unsigned(195, 10) ) ELSE
                     delay_pipeline(230) WHEN ( cur_count = to_unsigned(196, 10) ) ELSE
                     delay_pipeline(231) WHEN ( cur_count = to_unsigned(197, 10) ) ELSE
                     delay_pipeline(232) WHEN ( cur_count = to_unsigned(198, 10) ) ELSE
                     delay_pipeline(233) WHEN ( cur_count = to_unsigned(199, 10) ) ELSE
                     delay_pipeline(234) WHEN ( cur_count = to_unsigned(200, 10) ) ELSE
                     delay_pipeline(235) WHEN ( cur_count = to_unsigned(201, 10) ) ELSE
                     delay_pipeline(236) WHEN ( cur_count = to_unsigned(202, 10) ) ELSE
                     delay_pipeline(237) WHEN ( cur_count = to_unsigned(203, 10) ) ELSE
                     delay_pipeline(238) WHEN ( cur_count = to_unsigned(204, 10) ) ELSE
                     delay_pipeline(239) WHEN ( cur_count = to_unsigned(205, 10) ) ELSE
                     delay_pipeline(240) WHEN ( cur_count = to_unsigned(206, 10) ) ELSE
                     delay_pipeline(241) WHEN ( cur_count = to_unsigned(207, 10) ) ELSE
                     delay_pipeline(242) WHEN ( cur_count = to_unsigned(208, 10) ) ELSE
                     delay_pipeline(243) WHEN ( cur_count = to_unsigned(209, 10) ) ELSE
                     delay_pipeline(244) WHEN ( cur_count = to_unsigned(210, 10) ) ELSE
                     delay_pipeline(245) WHEN ( cur_count = to_unsigned(211, 10) ) ELSE
                     delay_pipeline(246) WHEN ( cur_count = to_unsigned(212, 10) ) ELSE
                     delay_pipeline(247) WHEN ( cur_count = to_unsigned(213, 10) ) ELSE
                     delay_pipeline(248) WHEN ( cur_count = to_unsigned(214, 10) ) ELSE
                     delay_pipeline(249) WHEN ( cur_count = to_unsigned(215, 10) ) ELSE
                     delay_pipeline(251) WHEN ( cur_count = to_unsigned(216, 10) ) ELSE
                     delay_pipeline(252) WHEN ( cur_count = to_unsigned(217, 10) ) ELSE
                     delay_pipeline(253) WHEN ( cur_count = to_unsigned(218, 10) ) ELSE
                     delay_pipeline(254) WHEN ( cur_count = to_unsigned(219, 10) ) ELSE
                     delay_pipeline(255) WHEN ( cur_count = to_unsigned(220, 10) ) ELSE
                     delay_pipeline(256) WHEN ( cur_count = to_unsigned(221, 10) ) ELSE
                     delay_pipeline(257) WHEN ( cur_count = to_unsigned(222, 10) ) ELSE
                     delay_pipeline(258) WHEN ( cur_count = to_unsigned(223, 10) ) ELSE
                     delay_pipeline(259) WHEN ( cur_count = to_unsigned(224, 10) ) ELSE
                     delay_pipeline(260) WHEN ( cur_count = to_unsigned(225, 10) ) ELSE
                     delay_pipeline(261) WHEN ( cur_count = to_unsigned(226, 10) ) ELSE
                     delay_pipeline(262) WHEN ( cur_count = to_unsigned(227, 10) ) ELSE
                     delay_pipeline(263) WHEN ( cur_count = to_unsigned(228, 10) ) ELSE
                     delay_pipeline(264) WHEN ( cur_count = to_unsigned(229, 10) ) ELSE
                     delay_pipeline(265) WHEN ( cur_count = to_unsigned(230, 10) ) ELSE
                     delay_pipeline(266) WHEN ( cur_count = to_unsigned(231, 10) ) ELSE
                     delay_pipeline(267) WHEN ( cur_count = to_unsigned(232, 10) ) ELSE
                     delay_pipeline(268) WHEN ( cur_count = to_unsigned(233, 10) ) ELSE
                     delay_pipeline(269) WHEN ( cur_count = to_unsigned(234, 10) ) ELSE
                     delay_pipeline(270) WHEN ( cur_count = to_unsigned(235, 10) ) ELSE
                     delay_pipeline(271) WHEN ( cur_count = to_unsigned(236, 10) ) ELSE
                     delay_pipeline(272) WHEN ( cur_count = to_unsigned(237, 10) ) ELSE
                     delay_pipeline(273) WHEN ( cur_count = to_unsigned(238, 10) ) ELSE
                     delay_pipeline(274) WHEN ( cur_count = to_unsigned(239, 10) ) ELSE
                     delay_pipeline(275) WHEN ( cur_count = to_unsigned(240, 10) ) ELSE
                     delay_pipeline(276) WHEN ( cur_count = to_unsigned(241, 10) ) ELSE
                     delay_pipeline(277) WHEN ( cur_count = to_unsigned(242, 10) ) ELSE
                     delay_pipeline(278) WHEN ( cur_count = to_unsigned(243, 10) ) ELSE
                     delay_pipeline(279) WHEN ( cur_count = to_unsigned(244, 10) ) ELSE
                     delay_pipeline(280) WHEN ( cur_count = to_unsigned(245, 10) ) ELSE
                     delay_pipeline(281) WHEN ( cur_count = to_unsigned(246, 10) ) ELSE
                     delay_pipeline(282) WHEN ( cur_count = to_unsigned(247, 10) ) ELSE
                     delay_pipeline(283) WHEN ( cur_count = to_unsigned(248, 10) ) ELSE
                     delay_pipeline(284) WHEN ( cur_count = to_unsigned(249, 10) ) ELSE
                     delay_pipeline(285) WHEN ( cur_count = to_unsigned(250, 10) ) ELSE
                     delay_pipeline(286) WHEN ( cur_count = to_unsigned(251, 10) ) ELSE
                     delay_pipeline(287) WHEN ( cur_count = to_unsigned(252, 10) ) ELSE
                     delay_pipeline(288) WHEN ( cur_count = to_unsigned(253, 10) ) ELSE
                     delay_pipeline(289) WHEN ( cur_count = to_unsigned(254, 10) ) ELSE
                     delay_pipeline(290) WHEN ( cur_count = to_unsigned(255, 10) ) ELSE
                     delay_pipeline(291) WHEN ( cur_count = to_unsigned(256, 10) ) ELSE
                     delay_pipeline(292) WHEN ( cur_count = to_unsigned(257, 10) ) ELSE
                     delay_pipeline(293) WHEN ( cur_count = to_unsigned(258, 10) ) ELSE
                     delay_pipeline(294) WHEN ( cur_count = to_unsigned(259, 10) ) ELSE
                     delay_pipeline(295) WHEN ( cur_count = to_unsigned(260, 10) ) ELSE
                     delay_pipeline(296) WHEN ( cur_count = to_unsigned(261, 10) ) ELSE
                     delay_pipeline(297) WHEN ( cur_count = to_unsigned(262, 10) ) ELSE
                     delay_pipeline(299) WHEN ( cur_count = to_unsigned(263, 10) ) ELSE
                     delay_pipeline(300) WHEN ( cur_count = to_unsigned(264, 10) ) ELSE
                     delay_pipeline(301) WHEN ( cur_count = to_unsigned(265, 10) ) ELSE
                     delay_pipeline(302) WHEN ( cur_count = to_unsigned(266, 10) ) ELSE
                     delay_pipeline(303) WHEN ( cur_count = to_unsigned(267, 10) ) ELSE
                     delay_pipeline(304) WHEN ( cur_count = to_unsigned(268, 10) ) ELSE
                     delay_pipeline(305) WHEN ( cur_count = to_unsigned(269, 10) ) ELSE
                     delay_pipeline(306) WHEN ( cur_count = to_unsigned(270, 10) ) ELSE
                     delay_pipeline(307) WHEN ( cur_count = to_unsigned(271, 10) ) ELSE
                     delay_pipeline(308) WHEN ( cur_count = to_unsigned(272, 10) ) ELSE
                     delay_pipeline(309) WHEN ( cur_count = to_unsigned(273, 10) ) ELSE
                     delay_pipeline(310) WHEN ( cur_count = to_unsigned(274, 10) ) ELSE
                     delay_pipeline(311) WHEN ( cur_count = to_unsigned(275, 10) ) ELSE
                     delay_pipeline(312) WHEN ( cur_count = to_unsigned(276, 10) ) ELSE
                     delay_pipeline(313) WHEN ( cur_count = to_unsigned(277, 10) ) ELSE
                     delay_pipeline(314) WHEN ( cur_count = to_unsigned(278, 10) ) ELSE
                     delay_pipeline(315) WHEN ( cur_count = to_unsigned(279, 10) ) ELSE
                     delay_pipeline(316) WHEN ( cur_count = to_unsigned(280, 10) ) ELSE
                     delay_pipeline(317) WHEN ( cur_count = to_unsigned(281, 10) ) ELSE
                     delay_pipeline(318) WHEN ( cur_count = to_unsigned(282, 10) ) ELSE
                     delay_pipeline(319) WHEN ( cur_count = to_unsigned(283, 10) ) ELSE
                     delay_pipeline(320) WHEN ( cur_count = to_unsigned(284, 10) ) ELSE
                     delay_pipeline(321) WHEN ( cur_count = to_unsigned(285, 10) ) ELSE
                     delay_pipeline(322) WHEN ( cur_count = to_unsigned(286, 10) ) ELSE
                     delay_pipeline(323) WHEN ( cur_count = to_unsigned(287, 10) ) ELSE
                     delay_pipeline(324) WHEN ( cur_count = to_unsigned(288, 10) ) ELSE
                     delay_pipeline(325) WHEN ( cur_count = to_unsigned(289, 10) ) ELSE
                     delay_pipeline(326) WHEN ( cur_count = to_unsigned(290, 10) ) ELSE
                     delay_pipeline(327) WHEN ( cur_count = to_unsigned(291, 10) ) ELSE
                     delay_pipeline(328) WHEN ( cur_count = to_unsigned(292, 10) ) ELSE
                     delay_pipeline(329) WHEN ( cur_count = to_unsigned(293, 10) ) ELSE
                     delay_pipeline(330) WHEN ( cur_count = to_unsigned(294, 10) ) ELSE
                     delay_pipeline(331) WHEN ( cur_count = to_unsigned(295, 10) ) ELSE
                     delay_pipeline(332) WHEN ( cur_count = to_unsigned(296, 10) ) ELSE
                     delay_pipeline(333) WHEN ( cur_count = to_unsigned(297, 10) ) ELSE
                     delay_pipeline(334) WHEN ( cur_count = to_unsigned(298, 10) ) ELSE
                     delay_pipeline(335) WHEN ( cur_count = to_unsigned(299, 10) ) ELSE
                     delay_pipeline(336) WHEN ( cur_count = to_unsigned(300, 10) ) ELSE
                     delay_pipeline(337) WHEN ( cur_count = to_unsigned(301, 10) ) ELSE
                     delay_pipeline(338) WHEN ( cur_count = to_unsigned(302, 10) ) ELSE
                     delay_pipeline(339) WHEN ( cur_count = to_unsigned(303, 10) ) ELSE
                     delay_pipeline(340) WHEN ( cur_count = to_unsigned(304, 10) ) ELSE
                     delay_pipeline(341) WHEN ( cur_count = to_unsigned(305, 10) ) ELSE
                     delay_pipeline(342) WHEN ( cur_count = to_unsigned(306, 10) ) ELSE
                     delay_pipeline(343) WHEN ( cur_count = to_unsigned(307, 10) ) ELSE
                     delay_pipeline(344) WHEN ( cur_count = to_unsigned(308, 10) ) ELSE
                     delay_pipeline(345) WHEN ( cur_count = to_unsigned(309, 10) ) ELSE
                     delay_pipeline(346) WHEN ( cur_count = to_unsigned(310, 10) ) ELSE
                     delay_pipeline(347) WHEN ( cur_count = to_unsigned(311, 10) ) ELSE
                     delay_pipeline(348) WHEN ( cur_count = to_unsigned(312, 10) ) ELSE
                     delay_pipeline(349) WHEN ( cur_count = to_unsigned(313, 10) ) ELSE
                     delay_pipeline(350) WHEN ( cur_count = to_unsigned(314, 10) ) ELSE
                     delay_pipeline(351) WHEN ( cur_count = to_unsigned(315, 10) ) ELSE
                     delay_pipeline(352) WHEN ( cur_count = to_unsigned(316, 10) ) ELSE
                     delay_pipeline(353) WHEN ( cur_count = to_unsigned(317, 10) ) ELSE
                     delay_pipeline(354) WHEN ( cur_count = to_unsigned(318, 10) ) ELSE
                     delay_pipeline(355) WHEN ( cur_count = to_unsigned(319, 10) ) ELSE
                     delay_pipeline(356) WHEN ( cur_count = to_unsigned(320, 10) ) ELSE
                     delay_pipeline(357) WHEN ( cur_count = to_unsigned(321, 10) ) ELSE
                     delay_pipeline(358) WHEN ( cur_count = to_unsigned(322, 10) ) ELSE
                     delay_pipeline(359) WHEN ( cur_count = to_unsigned(323, 10) ) ELSE
                     delay_pipeline(360) WHEN ( cur_count = to_unsigned(324, 10) ) ELSE
                     delay_pipeline(361) WHEN ( cur_count = to_unsigned(325, 10) ) ELSE
                     delay_pipeline(362) WHEN ( cur_count = to_unsigned(326, 10) ) ELSE
                     delay_pipeline(363) WHEN ( cur_count = to_unsigned(327, 10) ) ELSE
                     delay_pipeline(364) WHEN ( cur_count = to_unsigned(328, 10) ) ELSE
                     delay_pipeline(365) WHEN ( cur_count = to_unsigned(329, 10) ) ELSE
                     delay_pipeline(366) WHEN ( cur_count = to_unsigned(330, 10) ) ELSE
                     delay_pipeline(367) WHEN ( cur_count = to_unsigned(331, 10) ) ELSE
                     delay_pipeline(368) WHEN ( cur_count = to_unsigned(332, 10) ) ELSE
                     delay_pipeline(369) WHEN ( cur_count = to_unsigned(333, 10) ) ELSE
                     delay_pipeline(370) WHEN ( cur_count = to_unsigned(334, 10) ) ELSE
                     delay_pipeline(371) WHEN ( cur_count = to_unsigned(335, 10) ) ELSE
                     delay_pipeline(372) WHEN ( cur_count = to_unsigned(336, 10) ) ELSE
                     delay_pipeline(373) WHEN ( cur_count = to_unsigned(337, 10) ) ELSE
                     delay_pipeline(374) WHEN ( cur_count = to_unsigned(338, 10) ) ELSE
                     delay_pipeline(375) WHEN ( cur_count = to_unsigned(339, 10) ) ELSE
                     delay_pipeline(376) WHEN ( cur_count = to_unsigned(340, 10) ) ELSE
                     delay_pipeline(377) WHEN ( cur_count = to_unsigned(341, 10) ) ELSE
                     delay_pipeline(378) WHEN ( cur_count = to_unsigned(342, 10) ) ELSE
                     delay_pipeline(379) WHEN ( cur_count = to_unsigned(343, 10) ) ELSE
                     delay_pipeline(380) WHEN ( cur_count = to_unsigned(344, 10) ) ELSE
                     delay_pipeline(381) WHEN ( cur_count = to_unsigned(345, 10) ) ELSE
                     delay_pipeline(382) WHEN ( cur_count = to_unsigned(346, 10) ) ELSE
                     delay_pipeline(383) WHEN ( cur_count = to_unsigned(347, 10) ) ELSE
                     delay_pipeline(384) WHEN ( cur_count = to_unsigned(348, 10) ) ELSE
                     delay_pipeline(385) WHEN ( cur_count = to_unsigned(349, 10) ) ELSE
                     delay_pipeline(386) WHEN ( cur_count = to_unsigned(350, 10) ) ELSE
                     delay_pipeline(387) WHEN ( cur_count = to_unsigned(351, 10) ) ELSE
                     delay_pipeline(388) WHEN ( cur_count = to_unsigned(352, 10) ) ELSE
                     delay_pipeline(389) WHEN ( cur_count = to_unsigned(353, 10) ) ELSE
                     delay_pipeline(390) WHEN ( cur_count = to_unsigned(354, 10) ) ELSE
                     delay_pipeline(391) WHEN ( cur_count = to_unsigned(355, 10) ) ELSE
                     delay_pipeline(392) WHEN ( cur_count = to_unsigned(356, 10) ) ELSE
                     delay_pipeline(393) WHEN ( cur_count = to_unsigned(357, 10) ) ELSE
                     delay_pipeline(394) WHEN ( cur_count = to_unsigned(358, 10) ) ELSE
                     delay_pipeline(396) WHEN ( cur_count = to_unsigned(359, 10) ) ELSE
                     delay_pipeline(397) WHEN ( cur_count = to_unsigned(360, 10) ) ELSE
                     delay_pipeline(398) WHEN ( cur_count = to_unsigned(361, 10) ) ELSE
                     delay_pipeline(399) WHEN ( cur_count = to_unsigned(362, 10) ) ELSE
                     delay_pipeline(400) WHEN ( cur_count = to_unsigned(363, 10) ) ELSE
                     delay_pipeline(401) WHEN ( cur_count = to_unsigned(364, 10) ) ELSE
                     delay_pipeline(402) WHEN ( cur_count = to_unsigned(365, 10) ) ELSE
                     delay_pipeline(403) WHEN ( cur_count = to_unsigned(366, 10) ) ELSE
                     delay_pipeline(404) WHEN ( cur_count = to_unsigned(367, 10) ) ELSE
                     delay_pipeline(405) WHEN ( cur_count = to_unsigned(368, 10) ) ELSE
                     delay_pipeline(406) WHEN ( cur_count = to_unsigned(369, 10) ) ELSE
                     delay_pipeline(407) WHEN ( cur_count = to_unsigned(370, 10) ) ELSE
                     delay_pipeline(408) WHEN ( cur_count = to_unsigned(371, 10) ) ELSE
                     delay_pipeline(409) WHEN ( cur_count = to_unsigned(372, 10) ) ELSE
                     delay_pipeline(410) WHEN ( cur_count = to_unsigned(373, 10) ) ELSE
                     delay_pipeline(411) WHEN ( cur_count = to_unsigned(374, 10) ) ELSE
                     delay_pipeline(412) WHEN ( cur_count = to_unsigned(375, 10) ) ELSE
                     delay_pipeline(413) WHEN ( cur_count = to_unsigned(376, 10) ) ELSE
                     delay_pipeline(414) WHEN ( cur_count = to_unsigned(377, 10) ) ELSE
                     delay_pipeline(415) WHEN ( cur_count = to_unsigned(378, 10) ) ELSE
                     delay_pipeline(416) WHEN ( cur_count = to_unsigned(379, 10) ) ELSE
                     delay_pipeline(417) WHEN ( cur_count = to_unsigned(380, 10) ) ELSE
                     delay_pipeline(418) WHEN ( cur_count = to_unsigned(381, 10) ) ELSE
                     delay_pipeline(419) WHEN ( cur_count = to_unsigned(382, 10) ) ELSE
                     delay_pipeline(420) WHEN ( cur_count = to_unsigned(383, 10) ) ELSE
                     delay_pipeline(421) WHEN ( cur_count = to_unsigned(384, 10) ) ELSE
                     delay_pipeline(422) WHEN ( cur_count = to_unsigned(385, 10) ) ELSE
                     delay_pipeline(423) WHEN ( cur_count = to_unsigned(386, 10) ) ELSE
                     delay_pipeline(424) WHEN ( cur_count = to_unsigned(387, 10) ) ELSE
                     delay_pipeline(425) WHEN ( cur_count = to_unsigned(388, 10) ) ELSE
                     delay_pipeline(426) WHEN ( cur_count = to_unsigned(389, 10) ) ELSE
                     delay_pipeline(427) WHEN ( cur_count = to_unsigned(390, 10) ) ELSE
                     delay_pipeline(428) WHEN ( cur_count = to_unsigned(391, 10) ) ELSE
                     delay_pipeline(429) WHEN ( cur_count = to_unsigned(392, 10) ) ELSE
                     delay_pipeline(430) WHEN ( cur_count = to_unsigned(393, 10) ) ELSE
                     delay_pipeline(431) WHEN ( cur_count = to_unsigned(394, 10) ) ELSE
                     delay_pipeline(432) WHEN ( cur_count = to_unsigned(395, 10) ) ELSE
                     delay_pipeline(433) WHEN ( cur_count = to_unsigned(396, 10) ) ELSE
                     delay_pipeline(434) WHEN ( cur_count = to_unsigned(397, 10) ) ELSE
                     delay_pipeline(435) WHEN ( cur_count = to_unsigned(398, 10) ) ELSE
                     delay_pipeline(436) WHEN ( cur_count = to_unsigned(399, 10) ) ELSE
                     delay_pipeline(437) WHEN ( cur_count = to_unsigned(400, 10) ) ELSE
                     delay_pipeline(438) WHEN ( cur_count = to_unsigned(401, 10) ) ELSE
                     delay_pipeline(439) WHEN ( cur_count = to_unsigned(402, 10) ) ELSE
                     delay_pipeline(440) WHEN ( cur_count = to_unsigned(403, 10) ) ELSE
                     delay_pipeline(441) WHEN ( cur_count = to_unsigned(404, 10) ) ELSE
                     delay_pipeline(442) WHEN ( cur_count = to_unsigned(405, 10) ) ELSE
                     delay_pipeline(444) WHEN ( cur_count = to_unsigned(406, 10) ) ELSE
                     delay_pipeline(445) WHEN ( cur_count = to_unsigned(407, 10) ) ELSE
                     delay_pipeline(446) WHEN ( cur_count = to_unsigned(408, 10) ) ELSE
                     delay_pipeline(447) WHEN ( cur_count = to_unsigned(409, 10) ) ELSE
                     delay_pipeline(448) WHEN ( cur_count = to_unsigned(410, 10) ) ELSE
                     delay_pipeline(449) WHEN ( cur_count = to_unsigned(411, 10) ) ELSE
                     delay_pipeline(450) WHEN ( cur_count = to_unsigned(412, 10) ) ELSE
                     delay_pipeline(451) WHEN ( cur_count = to_unsigned(413, 10) ) ELSE
                     delay_pipeline(452) WHEN ( cur_count = to_unsigned(414, 10) ) ELSE
                     delay_pipeline(453) WHEN ( cur_count = to_unsigned(415, 10) ) ELSE
                     delay_pipeline(454) WHEN ( cur_count = to_unsigned(416, 10) ) ELSE
                     delay_pipeline(455) WHEN ( cur_count = to_unsigned(417, 10) ) ELSE
                     delay_pipeline(456) WHEN ( cur_count = to_unsigned(418, 10) ) ELSE
                     delay_pipeline(457) WHEN ( cur_count = to_unsigned(419, 10) ) ELSE
                     delay_pipeline(458) WHEN ( cur_count = to_unsigned(420, 10) ) ELSE
                     delay_pipeline(459) WHEN ( cur_count = to_unsigned(421, 10) ) ELSE
                     delay_pipeline(460) WHEN ( cur_count = to_unsigned(422, 10) ) ELSE
                     delay_pipeline(461) WHEN ( cur_count = to_unsigned(423, 10) ) ELSE
                     delay_pipeline(462) WHEN ( cur_count = to_unsigned(424, 10) ) ELSE
                     delay_pipeline(463) WHEN ( cur_count = to_unsigned(425, 10) ) ELSE
                     delay_pipeline(464) WHEN ( cur_count = to_unsigned(426, 10) ) ELSE
                     delay_pipeline(465) WHEN ( cur_count = to_unsigned(427, 10) ) ELSE
                     delay_pipeline(466) WHEN ( cur_count = to_unsigned(428, 10) ) ELSE
                     delay_pipeline(467) WHEN ( cur_count = to_unsigned(429, 10) ) ELSE
                     delay_pipeline(468) WHEN ( cur_count = to_unsigned(430, 10) ) ELSE
                     delay_pipeline(469) WHEN ( cur_count = to_unsigned(431, 10) ) ELSE
                     delay_pipeline(470) WHEN ( cur_count = to_unsigned(432, 10) ) ELSE
                     delay_pipeline(471) WHEN ( cur_count = to_unsigned(433, 10) ) ELSE
                     delay_pipeline(472) WHEN ( cur_count = to_unsigned(434, 10) ) ELSE
                     delay_pipeline(473) WHEN ( cur_count = to_unsigned(435, 10) ) ELSE
                     delay_pipeline(474) WHEN ( cur_count = to_unsigned(436, 10) ) ELSE
                     delay_pipeline(475) WHEN ( cur_count = to_unsigned(437, 10) ) ELSE
                     delay_pipeline(476) WHEN ( cur_count = to_unsigned(438, 10) ) ELSE
                     delay_pipeline(477) WHEN ( cur_count = to_unsigned(439, 10) ) ELSE
                     delay_pipeline(478) WHEN ( cur_count = to_unsigned(440, 10) ) ELSE
                     delay_pipeline(479) WHEN ( cur_count = to_unsigned(441, 10) ) ELSE
                     delay_pipeline(480) WHEN ( cur_count = to_unsigned(442, 10) ) ELSE
                     delay_pipeline(481) WHEN ( cur_count = to_unsigned(443, 10) ) ELSE
                     delay_pipeline(482) WHEN ( cur_count = to_unsigned(444, 10) ) ELSE
                     delay_pipeline(483) WHEN ( cur_count = to_unsigned(445, 10) ) ELSE
                     delay_pipeline(484) WHEN ( cur_count = to_unsigned(446, 10) ) ELSE
                     delay_pipeline(485) WHEN ( cur_count = to_unsigned(447, 10) ) ELSE
                     delay_pipeline(486) WHEN ( cur_count = to_unsigned(448, 10) ) ELSE
                     delay_pipeline(487) WHEN ( cur_count = to_unsigned(449, 10) ) ELSE
                     delay_pipeline(488) WHEN ( cur_count = to_unsigned(450, 10) ) ELSE
                     delay_pipeline(489) WHEN ( cur_count = to_unsigned(451, 10) ) ELSE
                     delay_pipeline(490) WHEN ( cur_count = to_unsigned(452, 10) ) ELSE
                     delay_pipeline(493) WHEN ( cur_count = to_unsigned(453, 10) ) ELSE
                     delay_pipeline(494) WHEN ( cur_count = to_unsigned(454, 10) ) ELSE
                     delay_pipeline(495) WHEN ( cur_count = to_unsigned(455, 10) ) ELSE
                     delay_pipeline(496) WHEN ( cur_count = to_unsigned(456, 10) ) ELSE
                     delay_pipeline(497) WHEN ( cur_count = to_unsigned(457, 10) ) ELSE
                     delay_pipeline(498) WHEN ( cur_count = to_unsigned(458, 10) ) ELSE
                     delay_pipeline(499) WHEN ( cur_count = to_unsigned(459, 10) ) ELSE
                     delay_pipeline(500) WHEN ( cur_count = to_unsigned(460, 10) ) ELSE
                     delay_pipeline(501) WHEN ( cur_count = to_unsigned(461, 10) ) ELSE
                     delay_pipeline(502) WHEN ( cur_count = to_unsigned(462, 10) ) ELSE
                     delay_pipeline(503) WHEN ( cur_count = to_unsigned(463, 10) ) ELSE
                     delay_pipeline(504) WHEN ( cur_count = to_unsigned(464, 10) ) ELSE
                     delay_pipeline(505) WHEN ( cur_count = to_unsigned(465, 10) ) ELSE
                     delay_pipeline(506) WHEN ( cur_count = to_unsigned(466, 10) ) ELSE
                     delay_pipeline(507) WHEN ( cur_count = to_unsigned(467, 10) ) ELSE
                     delay_pipeline(508) WHEN ( cur_count = to_unsigned(468, 10) ) ELSE
                     delay_pipeline(509) WHEN ( cur_count = to_unsigned(469, 10) ) ELSE
                     delay_pipeline(510) WHEN ( cur_count = to_unsigned(470, 10) ) ELSE
                     delay_pipeline(511) WHEN ( cur_count = to_unsigned(471, 10) ) ELSE
                     delay_pipeline(512) WHEN ( cur_count = to_unsigned(472, 10) ) ELSE
                     delay_pipeline(513) WHEN ( cur_count = to_unsigned(473, 10) ) ELSE
                     delay_pipeline(514) WHEN ( cur_count = to_unsigned(474, 10) ) ELSE
                     delay_pipeline(515) WHEN ( cur_count = to_unsigned(475, 10) ) ELSE
                     delay_pipeline(516) WHEN ( cur_count = to_unsigned(476, 10) ) ELSE
                     delay_pipeline(517) WHEN ( cur_count = to_unsigned(477, 10) ) ELSE
                     delay_pipeline(518) WHEN ( cur_count = to_unsigned(478, 10) ) ELSE
                     delay_pipeline(519) WHEN ( cur_count = to_unsigned(479, 10) ) ELSE
                     delay_pipeline(520) WHEN ( cur_count = to_unsigned(480, 10) ) ELSE
                     delay_pipeline(521) WHEN ( cur_count = to_unsigned(481, 10) ) ELSE
                     delay_pipeline(522) WHEN ( cur_count = to_unsigned(482, 10) ) ELSE
                     delay_pipeline(523) WHEN ( cur_count = to_unsigned(483, 10) ) ELSE
                     delay_pipeline(524) WHEN ( cur_count = to_unsigned(484, 10) ) ELSE
                     delay_pipeline(525) WHEN ( cur_count = to_unsigned(485, 10) ) ELSE
                     delay_pipeline(526) WHEN ( cur_count = to_unsigned(486, 10) ) ELSE
                     delay_pipeline(527) WHEN ( cur_count = to_unsigned(487, 10) ) ELSE
                     delay_pipeline(528) WHEN ( cur_count = to_unsigned(488, 10) ) ELSE
                     delay_pipeline(529) WHEN ( cur_count = to_unsigned(489, 10) ) ELSE
                     delay_pipeline(530) WHEN ( cur_count = to_unsigned(490, 10) ) ELSE
                     delay_pipeline(531) WHEN ( cur_count = to_unsigned(491, 10) ) ELSE
                     delay_pipeline(532) WHEN ( cur_count = to_unsigned(492, 10) ) ELSE
                     delay_pipeline(533) WHEN ( cur_count = to_unsigned(493, 10) ) ELSE
                     delay_pipeline(534) WHEN ( cur_count = to_unsigned(494, 10) ) ELSE
                     delay_pipeline(535) WHEN ( cur_count = to_unsigned(495, 10) ) ELSE
                     delay_pipeline(536) WHEN ( cur_count = to_unsigned(496, 10) ) ELSE
                     delay_pipeline(537) WHEN ( cur_count = to_unsigned(497, 10) ) ELSE
                     delay_pipeline(542) WHEN ( cur_count = to_unsigned(498, 10) ) ELSE
                     delay_pipeline(543) WHEN ( cur_count = to_unsigned(499, 10) ) ELSE
                     delay_pipeline(544) WHEN ( cur_count = to_unsigned(500, 10) ) ELSE
                     delay_pipeline(545) WHEN ( cur_count = to_unsigned(501, 10) ) ELSE
                     delay_pipeline(546) WHEN ( cur_count = to_unsigned(502, 10) ) ELSE
                     delay_pipeline(547) WHEN ( cur_count = to_unsigned(503, 10) ) ELSE
                     delay_pipeline(548) WHEN ( cur_count = to_unsigned(504, 10) ) ELSE
                     delay_pipeline(549) WHEN ( cur_count = to_unsigned(505, 10) ) ELSE
                     delay_pipeline(550) WHEN ( cur_count = to_unsigned(506, 10) ) ELSE
                     delay_pipeline(551) WHEN ( cur_count = to_unsigned(507, 10) ) ELSE
                     delay_pipeline(552) WHEN ( cur_count = to_unsigned(508, 10) ) ELSE
                     delay_pipeline(553) WHEN ( cur_count = to_unsigned(509, 10) ) ELSE
                     delay_pipeline(554) WHEN ( cur_count = to_unsigned(510, 10) ) ELSE
                     delay_pipeline(555) WHEN ( cur_count = to_unsigned(511, 10) ) ELSE
                     delay_pipeline(556) WHEN ( cur_count = to_unsigned(512, 10) ) ELSE
                     delay_pipeline(557) WHEN ( cur_count = to_unsigned(513, 10) ) ELSE
                     delay_pipeline(558) WHEN ( cur_count = to_unsigned(514, 10) ) ELSE
                     delay_pipeline(559) WHEN ( cur_count = to_unsigned(515, 10) ) ELSE
                     delay_pipeline(560) WHEN ( cur_count = to_unsigned(516, 10) ) ELSE
                     delay_pipeline(561) WHEN ( cur_count = to_unsigned(517, 10) ) ELSE
                     delay_pipeline(562) WHEN ( cur_count = to_unsigned(518, 10) ) ELSE
                     delay_pipeline(563) WHEN ( cur_count = to_unsigned(519, 10) ) ELSE
                     delay_pipeline(564) WHEN ( cur_count = to_unsigned(520, 10) ) ELSE
                     delay_pipeline(565) WHEN ( cur_count = to_unsigned(521, 10) ) ELSE
                     delay_pipeline(566) WHEN ( cur_count = to_unsigned(522, 10) ) ELSE
                     delay_pipeline(567) WHEN ( cur_count = to_unsigned(523, 10) ) ELSE
                     delay_pipeline(568) WHEN ( cur_count = to_unsigned(524, 10) ) ELSE
                     delay_pipeline(569) WHEN ( cur_count = to_unsigned(525, 10) ) ELSE
                     delay_pipeline(570) WHEN ( cur_count = to_unsigned(526, 10) ) ELSE
                     delay_pipeline(571) WHEN ( cur_count = to_unsigned(527, 10) ) ELSE
                     delay_pipeline(572) WHEN ( cur_count = to_unsigned(528, 10) ) ELSE
                     delay_pipeline(573) WHEN ( cur_count = to_unsigned(529, 10) ) ELSE
                     delay_pipeline(574) WHEN ( cur_count = to_unsigned(530, 10) ) ELSE
                     delay_pipeline(575) WHEN ( cur_count = to_unsigned(531, 10) ) ELSE
                     delay_pipeline(576) WHEN ( cur_count = to_unsigned(532, 10) ) ELSE
                     delay_pipeline(577) WHEN ( cur_count = to_unsigned(533, 10) ) ELSE
                     delay_pipeline(578) WHEN ( cur_count = to_unsigned(534, 10) ) ELSE
                     delay_pipeline(579) WHEN ( cur_count = to_unsigned(535, 10) ) ELSE
                     delay_pipeline(580) WHEN ( cur_count = to_unsigned(536, 10) ) ELSE
                     delay_pipeline(581) WHEN ( cur_count = to_unsigned(537, 10) ) ELSE
                     delay_pipeline(582) WHEN ( cur_count = to_unsigned(538, 10) ) ELSE
                     delay_pipeline(583) WHEN ( cur_count = to_unsigned(539, 10) ) ELSE
                     delay_pipeline(591) WHEN ( cur_count = to_unsigned(540, 10) ) ELSE
                     delay_pipeline(592) WHEN ( cur_count = to_unsigned(541, 10) ) ELSE
                     delay_pipeline(593) WHEN ( cur_count = to_unsigned(542, 10) ) ELSE
                     delay_pipeline(594) WHEN ( cur_count = to_unsigned(543, 10) ) ELSE
                     delay_pipeline(595) WHEN ( cur_count = to_unsigned(544, 10) ) ELSE
                     delay_pipeline(596) WHEN ( cur_count = to_unsigned(545, 10) ) ELSE
                     delay_pipeline(597) WHEN ( cur_count = to_unsigned(546, 10) ) ELSE
                     delay_pipeline(598) WHEN ( cur_count = to_unsigned(547, 10) ) ELSE
                     delay_pipeline(599) WHEN ( cur_count = to_unsigned(548, 10) ) ELSE
                     delay_pipeline(600) WHEN ( cur_count = to_unsigned(549, 10) ) ELSE
                     delay_pipeline(601) WHEN ( cur_count = to_unsigned(550, 10) ) ELSE
                     delay_pipeline(602) WHEN ( cur_count = to_unsigned(551, 10) ) ELSE
                     delay_pipeline(603) WHEN ( cur_count = to_unsigned(552, 10) ) ELSE
                     delay_pipeline(604) WHEN ( cur_count = to_unsigned(553, 10) ) ELSE
                     delay_pipeline(605) WHEN ( cur_count = to_unsigned(554, 10) ) ELSE
                     delay_pipeline(606) WHEN ( cur_count = to_unsigned(555, 10) ) ELSE
                     delay_pipeline(607) WHEN ( cur_count = to_unsigned(556, 10) ) ELSE
                     delay_pipeline(608) WHEN ( cur_count = to_unsigned(557, 10) ) ELSE
                     delay_pipeline(609) WHEN ( cur_count = to_unsigned(558, 10) ) ELSE
                     delay_pipeline(610) WHEN ( cur_count = to_unsigned(559, 10) ) ELSE
                     delay_pipeline(611) WHEN ( cur_count = to_unsigned(560, 10) ) ELSE
                     delay_pipeline(612) WHEN ( cur_count = to_unsigned(561, 10) ) ELSE
                     delay_pipeline(613) WHEN ( cur_count = to_unsigned(562, 10) ) ELSE
                     delay_pipeline(614) WHEN ( cur_count = to_unsigned(563, 10) ) ELSE
                     delay_pipeline(615) WHEN ( cur_count = to_unsigned(564, 10) ) ELSE
                     delay_pipeline(616) WHEN ( cur_count = to_unsigned(565, 10) ) ELSE
                     delay_pipeline(617) WHEN ( cur_count = to_unsigned(566, 10) ) ELSE
                     delay_pipeline(618) WHEN ( cur_count = to_unsigned(567, 10) ) ELSE
                     delay_pipeline(619) WHEN ( cur_count = to_unsigned(568, 10) ) ELSE
                     delay_pipeline(620) WHEN ( cur_count = to_unsigned(569, 10) ) ELSE
                     delay_pipeline(621) WHEN ( cur_count = to_unsigned(570, 10) ) ELSE
                     delay_pipeline(622) WHEN ( cur_count = to_unsigned(571, 10) ) ELSE
                     delay_pipeline(623) WHEN ( cur_count = to_unsigned(572, 10) ) ELSE
                     delay_pipeline(624) WHEN ( cur_count = to_unsigned(573, 10) ) ELSE
                     delay_pipeline(625) WHEN ( cur_count = to_unsigned(574, 10) ) ELSE
                     delay_pipeline(626) WHEN ( cur_count = to_unsigned(575, 10) ) ELSE
                     delay_pipeline(627) WHEN ( cur_count = to_unsigned(576, 10) ) ELSE
                     delay_pipeline(628) WHEN ( cur_count = to_unsigned(577, 10) ) ELSE
                     delay_pipeline(642) WHEN ( cur_count = to_unsigned(578, 10) ) ELSE
                     delay_pipeline(643) WHEN ( cur_count = to_unsigned(579, 10) ) ELSE
                     delay_pipeline(644) WHEN ( cur_count = to_unsigned(580, 10) ) ELSE
                     delay_pipeline(645) WHEN ( cur_count = to_unsigned(581, 10) ) ELSE
                     delay_pipeline(646) WHEN ( cur_count = to_unsigned(582, 10) ) ELSE
                     delay_pipeline(647) WHEN ( cur_count = to_unsigned(583, 10) ) ELSE
                     delay_pipeline(648) WHEN ( cur_count = to_unsigned(584, 10) ) ELSE
                     delay_pipeline(649) WHEN ( cur_count = to_unsigned(585, 10) ) ELSE
                     delay_pipeline(650) WHEN ( cur_count = to_unsigned(586, 10) ) ELSE
                     delay_pipeline(651) WHEN ( cur_count = to_unsigned(587, 10) ) ELSE
                     delay_pipeline(652) WHEN ( cur_count = to_unsigned(588, 10) ) ELSE
                     delay_pipeline(653) WHEN ( cur_count = to_unsigned(589, 10) ) ELSE
                     delay_pipeline(654) WHEN ( cur_count = to_unsigned(590, 10) ) ELSE
                     delay_pipeline(655) WHEN ( cur_count = to_unsigned(591, 10) ) ELSE
                     delay_pipeline(656) WHEN ( cur_count = to_unsigned(592, 10) ) ELSE
                     delay_pipeline(657) WHEN ( cur_count = to_unsigned(593, 10) ) ELSE
                     delay_pipeline(658) WHEN ( cur_count = to_unsigned(594, 10) ) ELSE
                     delay_pipeline(659) WHEN ( cur_count = to_unsigned(595, 10) ) ELSE
                     delay_pipeline(660) WHEN ( cur_count = to_unsigned(596, 10) ) ELSE
                     delay_pipeline(661) WHEN ( cur_count = to_unsigned(597, 10) ) ELSE
                     delay_pipeline(662) WHEN ( cur_count = to_unsigned(598, 10) ) ELSE
                     delay_pipeline(663) WHEN ( cur_count = to_unsigned(599, 10) ) ELSE
                     delay_pipeline(664) WHEN ( cur_count = to_unsigned(600, 10) ) ELSE
                     delay_pipeline(665) WHEN ( cur_count = to_unsigned(601, 10) ) ELSE
                     delay_pipeline(666) WHEN ( cur_count = to_unsigned(602, 10) ) ELSE
                     delay_pipeline(667) WHEN ( cur_count = to_unsigned(603, 10) ) ELSE
                     delay_pipeline(668) WHEN ( cur_count = to_unsigned(604, 10) ) ELSE
                     delay_pipeline(669) WHEN ( cur_count = to_unsigned(605, 10) ) ELSE
                     delay_pipeline(670) WHEN ( cur_count = to_unsigned(606, 10) ) ELSE
                     delay_pipeline(671) WHEN ( cur_count = to_unsigned(607, 10) ) ELSE
                     delay_pipeline(672) WHEN ( cur_count = to_unsigned(608, 10) ) ELSE
                     delay_pipeline(673) WHEN ( cur_count = to_unsigned(609, 10) ) ELSE
                     delay_pipeline(674) WHEN ( cur_count = to_unsigned(610, 10) ) ELSE
                     delay_pipeline(675) WHEN ( cur_count = to_unsigned(611, 10) ) ELSE
                     delay_pipeline(676) WHEN ( cur_count = to_unsigned(612, 10) ) ELSE
                     delay_pipeline(685) WHEN ( cur_count = to_unsigned(613, 10) ) ELSE
                     delay_pipeline(686) WHEN ( cur_count = to_unsigned(614, 10) ) ELSE
                     delay_pipeline(687) WHEN ( cur_count = to_unsigned(615, 10) ) ELSE
                     delay_pipeline(688) WHEN ( cur_count = to_unsigned(616, 10) ) ELSE
                     delay_pipeline(689) WHEN ( cur_count = to_unsigned(617, 10) ) ELSE
                     delay_pipeline(690) WHEN ( cur_count = to_unsigned(618, 10) ) ELSE
                     delay_pipeline(691) WHEN ( cur_count = to_unsigned(619, 10) ) ELSE
                     delay_pipeline(692) WHEN ( cur_count = to_unsigned(620, 10) ) ELSE
                     delay_pipeline(693);

  --   ------------------ Serial partition # 1 ------------------

  product_1_mux <= coeff1 WHEN ( cur_count = to_unsigned(0, 10) ) ELSE
                        coeff2 WHEN ( cur_count = to_unsigned(1, 10) ) ELSE
                        coeff3 WHEN ( cur_count = to_unsigned(2, 10) ) ELSE
                        coeff4 WHEN ( cur_count = to_unsigned(3, 10) ) ELSE
                        coeff5 WHEN ( cur_count = to_unsigned(4, 10) ) ELSE
                        coeff6 WHEN ( cur_count = to_unsigned(5, 10) ) ELSE
                        coeff7 WHEN ( cur_count = to_unsigned(6, 10) ) ELSE
                        coeff8 WHEN ( cur_count = to_unsigned(7, 10) ) ELSE
                        coeff9 WHEN ( cur_count = to_unsigned(8, 10) ) ELSE
                        coeff18 WHEN ( cur_count = to_unsigned(9, 10) ) ELSE
                        coeff19 WHEN ( cur_count = to_unsigned(10, 10) ) ELSE
                        coeff20 WHEN ( cur_count = to_unsigned(11, 10) ) ELSE
                        coeff21 WHEN ( cur_count = to_unsigned(12, 10) ) ELSE
                        coeff22 WHEN ( cur_count = to_unsigned(13, 10) ) ELSE
                        coeff23 WHEN ( cur_count = to_unsigned(14, 10) ) ELSE
                        coeff24 WHEN ( cur_count = to_unsigned(15, 10) ) ELSE
                        coeff25 WHEN ( cur_count = to_unsigned(16, 10) ) ELSE
                        coeff26 WHEN ( cur_count = to_unsigned(17, 10) ) ELSE
                        coeff27 WHEN ( cur_count = to_unsigned(18, 10) ) ELSE
                        coeff28 WHEN ( cur_count = to_unsigned(19, 10) ) ELSE
                        coeff29 WHEN ( cur_count = to_unsigned(20, 10) ) ELSE
                        coeff30 WHEN ( cur_count = to_unsigned(21, 10) ) ELSE
                        coeff31 WHEN ( cur_count = to_unsigned(22, 10) ) ELSE
                        coeff32 WHEN ( cur_count = to_unsigned(23, 10) ) ELSE
                        coeff33 WHEN ( cur_count = to_unsigned(24, 10) ) ELSE
                        coeff34 WHEN ( cur_count = to_unsigned(25, 10) ) ELSE
                        coeff35 WHEN ( cur_count = to_unsigned(26, 10) ) ELSE
                        coeff36 WHEN ( cur_count = to_unsigned(27, 10) ) ELSE
                        coeff37 WHEN ( cur_count = to_unsigned(28, 10) ) ELSE
                        coeff38 WHEN ( cur_count = to_unsigned(29, 10) ) ELSE
                        coeff39 WHEN ( cur_count = to_unsigned(30, 10) ) ELSE
                        coeff40 WHEN ( cur_count = to_unsigned(31, 10) ) ELSE
                        coeff41 WHEN ( cur_count = to_unsigned(32, 10) ) ELSE
                        coeff42 WHEN ( cur_count = to_unsigned(33, 10) ) ELSE
                        coeff43 WHEN ( cur_count = to_unsigned(34, 10) ) ELSE
                        coeff44 WHEN ( cur_count = to_unsigned(35, 10) ) ELSE
                        coeff45 WHEN ( cur_count = to_unsigned(36, 10) ) ELSE
                        coeff46 WHEN ( cur_count = to_unsigned(37, 10) ) ELSE
                        coeff47 WHEN ( cur_count = to_unsigned(38, 10) ) ELSE
                        coeff48 WHEN ( cur_count = to_unsigned(39, 10) ) ELSE
                        coeff49 WHEN ( cur_count = to_unsigned(40, 10) ) ELSE
                        coeff50 WHEN ( cur_count = to_unsigned(41, 10) ) ELSE
                        coeff51 WHEN ( cur_count = to_unsigned(42, 10) ) ELSE
                        coeff52 WHEN ( cur_count = to_unsigned(43, 10) ) ELSE
                        coeff66 WHEN ( cur_count = to_unsigned(44, 10) ) ELSE
                        coeff67 WHEN ( cur_count = to_unsigned(45, 10) ) ELSE
                        coeff68 WHEN ( cur_count = to_unsigned(46, 10) ) ELSE
                        coeff69 WHEN ( cur_count = to_unsigned(47, 10) ) ELSE
                        coeff70 WHEN ( cur_count = to_unsigned(48, 10) ) ELSE
                        coeff71 WHEN ( cur_count = to_unsigned(49, 10) ) ELSE
                        coeff72 WHEN ( cur_count = to_unsigned(50, 10) ) ELSE
                        coeff73 WHEN ( cur_count = to_unsigned(51, 10) ) ELSE
                        coeff74 WHEN ( cur_count = to_unsigned(52, 10) ) ELSE
                        coeff75 WHEN ( cur_count = to_unsigned(53, 10) ) ELSE
                        coeff76 WHEN ( cur_count = to_unsigned(54, 10) ) ELSE
                        coeff77 WHEN ( cur_count = to_unsigned(55, 10) ) ELSE
                        coeff78 WHEN ( cur_count = to_unsigned(56, 10) ) ELSE
                        coeff79 WHEN ( cur_count = to_unsigned(57, 10) ) ELSE
                        coeff80 WHEN ( cur_count = to_unsigned(58, 10) ) ELSE
                        coeff81 WHEN ( cur_count = to_unsigned(59, 10) ) ELSE
                        coeff82 WHEN ( cur_count = to_unsigned(60, 10) ) ELSE
                        coeff83 WHEN ( cur_count = to_unsigned(61, 10) ) ELSE
                        coeff84 WHEN ( cur_count = to_unsigned(62, 10) ) ELSE
                        coeff85 WHEN ( cur_count = to_unsigned(63, 10) ) ELSE
                        coeff86 WHEN ( cur_count = to_unsigned(64, 10) ) ELSE
                        coeff87 WHEN ( cur_count = to_unsigned(65, 10) ) ELSE
                        coeff88 WHEN ( cur_count = to_unsigned(66, 10) ) ELSE
                        coeff89 WHEN ( cur_count = to_unsigned(67, 10) ) ELSE
                        coeff90 WHEN ( cur_count = to_unsigned(68, 10) ) ELSE
                        coeff91 WHEN ( cur_count = to_unsigned(69, 10) ) ELSE
                        coeff92 WHEN ( cur_count = to_unsigned(70, 10) ) ELSE
                        coeff93 WHEN ( cur_count = to_unsigned(71, 10) ) ELSE
                        coeff94 WHEN ( cur_count = to_unsigned(72, 10) ) ELSE
                        coeff95 WHEN ( cur_count = to_unsigned(73, 10) ) ELSE
                        coeff96 WHEN ( cur_count = to_unsigned(74, 10) ) ELSE
                        coeff97 WHEN ( cur_count = to_unsigned(75, 10) ) ELSE
                        coeff98 WHEN ( cur_count = to_unsigned(76, 10) ) ELSE
                        coeff99 WHEN ( cur_count = to_unsigned(77, 10) ) ELSE
                        coeff100 WHEN ( cur_count = to_unsigned(78, 10) ) ELSE
                        coeff101 WHEN ( cur_count = to_unsigned(79, 10) ) ELSE
                        coeff102 WHEN ( cur_count = to_unsigned(80, 10) ) ELSE
                        coeff103 WHEN ( cur_count = to_unsigned(81, 10) ) ELSE
                        coeff111 WHEN ( cur_count = to_unsigned(82, 10) ) ELSE
                        coeff112 WHEN ( cur_count = to_unsigned(83, 10) ) ELSE
                        coeff113 WHEN ( cur_count = to_unsigned(84, 10) ) ELSE
                        coeff114 WHEN ( cur_count = to_unsigned(85, 10) ) ELSE
                        coeff115 WHEN ( cur_count = to_unsigned(86, 10) ) ELSE
                        coeff116 WHEN ( cur_count = to_unsigned(87, 10) ) ELSE
                        coeff117 WHEN ( cur_count = to_unsigned(88, 10) ) ELSE
                        coeff118 WHEN ( cur_count = to_unsigned(89, 10) ) ELSE
                        coeff119 WHEN ( cur_count = to_unsigned(90, 10) ) ELSE
                        coeff120 WHEN ( cur_count = to_unsigned(91, 10) ) ELSE
                        coeff121 WHEN ( cur_count = to_unsigned(92, 10) ) ELSE
                        coeff122 WHEN ( cur_count = to_unsigned(93, 10) ) ELSE
                        coeff123 WHEN ( cur_count = to_unsigned(94, 10) ) ELSE
                        coeff124 WHEN ( cur_count = to_unsigned(95, 10) ) ELSE
                        coeff125 WHEN ( cur_count = to_unsigned(96, 10) ) ELSE
                        coeff126 WHEN ( cur_count = to_unsigned(97, 10) ) ELSE
                        coeff127 WHEN ( cur_count = to_unsigned(98, 10) ) ELSE
                        coeff128 WHEN ( cur_count = to_unsigned(99, 10) ) ELSE
                        coeff129 WHEN ( cur_count = to_unsigned(100, 10) ) ELSE
                        coeff130 WHEN ( cur_count = to_unsigned(101, 10) ) ELSE
                        coeff131 WHEN ( cur_count = to_unsigned(102, 10) ) ELSE
                        coeff132 WHEN ( cur_count = to_unsigned(103, 10) ) ELSE
                        coeff133 WHEN ( cur_count = to_unsigned(104, 10) ) ELSE
                        coeff134 WHEN ( cur_count = to_unsigned(105, 10) ) ELSE
                        coeff135 WHEN ( cur_count = to_unsigned(106, 10) ) ELSE
                        coeff136 WHEN ( cur_count = to_unsigned(107, 10) ) ELSE
                        coeff137 WHEN ( cur_count = to_unsigned(108, 10) ) ELSE
                        coeff138 WHEN ( cur_count = to_unsigned(109, 10) ) ELSE
                        coeff139 WHEN ( cur_count = to_unsigned(110, 10) ) ELSE
                        coeff140 WHEN ( cur_count = to_unsigned(111, 10) ) ELSE
                        coeff141 WHEN ( cur_count = to_unsigned(112, 10) ) ELSE
                        coeff142 WHEN ( cur_count = to_unsigned(113, 10) ) ELSE
                        coeff143 WHEN ( cur_count = to_unsigned(114, 10) ) ELSE
                        coeff144 WHEN ( cur_count = to_unsigned(115, 10) ) ELSE
                        coeff145 WHEN ( cur_count = to_unsigned(116, 10) ) ELSE
                        coeff146 WHEN ( cur_count = to_unsigned(117, 10) ) ELSE
                        coeff147 WHEN ( cur_count = to_unsigned(118, 10) ) ELSE
                        coeff148 WHEN ( cur_count = to_unsigned(119, 10) ) ELSE
                        coeff149 WHEN ( cur_count = to_unsigned(120, 10) ) ELSE
                        coeff150 WHEN ( cur_count = to_unsigned(121, 10) ) ELSE
                        coeff151 WHEN ( cur_count = to_unsigned(122, 10) ) ELSE
                        coeff152 WHEN ( cur_count = to_unsigned(123, 10) ) ELSE
                        coeff157 WHEN ( cur_count = to_unsigned(124, 10) ) ELSE
                        coeff158 WHEN ( cur_count = to_unsigned(125, 10) ) ELSE
                        coeff159 WHEN ( cur_count = to_unsigned(126, 10) ) ELSE
                        coeff160 WHEN ( cur_count = to_unsigned(127, 10) ) ELSE
                        coeff161 WHEN ( cur_count = to_unsigned(128, 10) ) ELSE
                        coeff162 WHEN ( cur_count = to_unsigned(129, 10) ) ELSE
                        coeff163 WHEN ( cur_count = to_unsigned(130, 10) ) ELSE
                        coeff164 WHEN ( cur_count = to_unsigned(131, 10) ) ELSE
                        coeff165 WHEN ( cur_count = to_unsigned(132, 10) ) ELSE
                        coeff166 WHEN ( cur_count = to_unsigned(133, 10) ) ELSE
                        coeff167 WHEN ( cur_count = to_unsigned(134, 10) ) ELSE
                        coeff168 WHEN ( cur_count = to_unsigned(135, 10) ) ELSE
                        coeff169 WHEN ( cur_count = to_unsigned(136, 10) ) ELSE
                        coeff170 WHEN ( cur_count = to_unsigned(137, 10) ) ELSE
                        coeff171 WHEN ( cur_count = to_unsigned(138, 10) ) ELSE
                        coeff172 WHEN ( cur_count = to_unsigned(139, 10) ) ELSE
                        coeff173 WHEN ( cur_count = to_unsigned(140, 10) ) ELSE
                        coeff174 WHEN ( cur_count = to_unsigned(141, 10) ) ELSE
                        coeff175 WHEN ( cur_count = to_unsigned(142, 10) ) ELSE
                        coeff176 WHEN ( cur_count = to_unsigned(143, 10) ) ELSE
                        coeff177 WHEN ( cur_count = to_unsigned(144, 10) ) ELSE
                        coeff178 WHEN ( cur_count = to_unsigned(145, 10) ) ELSE
                        coeff179 WHEN ( cur_count = to_unsigned(146, 10) ) ELSE
                        coeff180 WHEN ( cur_count = to_unsigned(147, 10) ) ELSE
                        coeff181 WHEN ( cur_count = to_unsigned(148, 10) ) ELSE
                        coeff182 WHEN ( cur_count = to_unsigned(149, 10) ) ELSE
                        coeff183 WHEN ( cur_count = to_unsigned(150, 10) ) ELSE
                        coeff184 WHEN ( cur_count = to_unsigned(151, 10) ) ELSE
                        coeff185 WHEN ( cur_count = to_unsigned(152, 10) ) ELSE
                        coeff186 WHEN ( cur_count = to_unsigned(153, 10) ) ELSE
                        coeff187 WHEN ( cur_count = to_unsigned(154, 10) ) ELSE
                        coeff188 WHEN ( cur_count = to_unsigned(155, 10) ) ELSE
                        coeff189 WHEN ( cur_count = to_unsigned(156, 10) ) ELSE
                        coeff190 WHEN ( cur_count = to_unsigned(157, 10) ) ELSE
                        coeff191 WHEN ( cur_count = to_unsigned(158, 10) ) ELSE
                        coeff192 WHEN ( cur_count = to_unsigned(159, 10) ) ELSE
                        coeff193 WHEN ( cur_count = to_unsigned(160, 10) ) ELSE
                        coeff194 WHEN ( cur_count = to_unsigned(161, 10) ) ELSE
                        coeff195 WHEN ( cur_count = to_unsigned(162, 10) ) ELSE
                        coeff196 WHEN ( cur_count = to_unsigned(163, 10) ) ELSE
                        coeff197 WHEN ( cur_count = to_unsigned(164, 10) ) ELSE
                        coeff198 WHEN ( cur_count = to_unsigned(165, 10) ) ELSE
                        coeff199 WHEN ( cur_count = to_unsigned(166, 10) ) ELSE
                        coeff200 WHEN ( cur_count = to_unsigned(167, 10) ) ELSE
                        coeff201 WHEN ( cur_count = to_unsigned(168, 10) ) ELSE
                        coeff204 WHEN ( cur_count = to_unsigned(169, 10) ) ELSE
                        coeff205 WHEN ( cur_count = to_unsigned(170, 10) ) ELSE
                        coeff206 WHEN ( cur_count = to_unsigned(171, 10) ) ELSE
                        coeff207 WHEN ( cur_count = to_unsigned(172, 10) ) ELSE
                        coeff208 WHEN ( cur_count = to_unsigned(173, 10) ) ELSE
                        coeff209 WHEN ( cur_count = to_unsigned(174, 10) ) ELSE
                        coeff210 WHEN ( cur_count = to_unsigned(175, 10) ) ELSE
                        coeff211 WHEN ( cur_count = to_unsigned(176, 10) ) ELSE
                        coeff212 WHEN ( cur_count = to_unsigned(177, 10) ) ELSE
                        coeff213 WHEN ( cur_count = to_unsigned(178, 10) ) ELSE
                        coeff214 WHEN ( cur_count = to_unsigned(179, 10) ) ELSE
                        coeff215 WHEN ( cur_count = to_unsigned(180, 10) ) ELSE
                        coeff216 WHEN ( cur_count = to_unsigned(181, 10) ) ELSE
                        coeff217 WHEN ( cur_count = to_unsigned(182, 10) ) ELSE
                        coeff218 WHEN ( cur_count = to_unsigned(183, 10) ) ELSE
                        coeff219 WHEN ( cur_count = to_unsigned(184, 10) ) ELSE
                        coeff220 WHEN ( cur_count = to_unsigned(185, 10) ) ELSE
                        coeff221 WHEN ( cur_count = to_unsigned(186, 10) ) ELSE
                        coeff222 WHEN ( cur_count = to_unsigned(187, 10) ) ELSE
                        coeff223 WHEN ( cur_count = to_unsigned(188, 10) ) ELSE
                        coeff224 WHEN ( cur_count = to_unsigned(189, 10) ) ELSE
                        coeff225 WHEN ( cur_count = to_unsigned(190, 10) ) ELSE
                        coeff226 WHEN ( cur_count = to_unsigned(191, 10) ) ELSE
                        coeff227 WHEN ( cur_count = to_unsigned(192, 10) ) ELSE
                        coeff228 WHEN ( cur_count = to_unsigned(193, 10) ) ELSE
                        coeff229 WHEN ( cur_count = to_unsigned(194, 10) ) ELSE
                        coeff230 WHEN ( cur_count = to_unsigned(195, 10) ) ELSE
                        coeff231 WHEN ( cur_count = to_unsigned(196, 10) ) ELSE
                        coeff232 WHEN ( cur_count = to_unsigned(197, 10) ) ELSE
                        coeff233 WHEN ( cur_count = to_unsigned(198, 10) ) ELSE
                        coeff234 WHEN ( cur_count = to_unsigned(199, 10) ) ELSE
                        coeff235 WHEN ( cur_count = to_unsigned(200, 10) ) ELSE
                        coeff236 WHEN ( cur_count = to_unsigned(201, 10) ) ELSE
                        coeff237 WHEN ( cur_count = to_unsigned(202, 10) ) ELSE
                        coeff238 WHEN ( cur_count = to_unsigned(203, 10) ) ELSE
                        coeff239 WHEN ( cur_count = to_unsigned(204, 10) ) ELSE
                        coeff240 WHEN ( cur_count = to_unsigned(205, 10) ) ELSE
                        coeff241 WHEN ( cur_count = to_unsigned(206, 10) ) ELSE
                        coeff242 WHEN ( cur_count = to_unsigned(207, 10) ) ELSE
                        coeff243 WHEN ( cur_count = to_unsigned(208, 10) ) ELSE
                        coeff244 WHEN ( cur_count = to_unsigned(209, 10) ) ELSE
                        coeff245 WHEN ( cur_count = to_unsigned(210, 10) ) ELSE
                        coeff246 WHEN ( cur_count = to_unsigned(211, 10) ) ELSE
                        coeff247 WHEN ( cur_count = to_unsigned(212, 10) ) ELSE
                        coeff248 WHEN ( cur_count = to_unsigned(213, 10) ) ELSE
                        coeff249 WHEN ( cur_count = to_unsigned(214, 10) ) ELSE
                        coeff250 WHEN ( cur_count = to_unsigned(215, 10) ) ELSE
                        coeff252 WHEN ( cur_count = to_unsigned(216, 10) ) ELSE
                        coeff253 WHEN ( cur_count = to_unsigned(217, 10) ) ELSE
                        coeff254 WHEN ( cur_count = to_unsigned(218, 10) ) ELSE
                        coeff255 WHEN ( cur_count = to_unsigned(219, 10) ) ELSE
                        coeff256 WHEN ( cur_count = to_unsigned(220, 10) ) ELSE
                        coeff257 WHEN ( cur_count = to_unsigned(221, 10) ) ELSE
                        coeff258 WHEN ( cur_count = to_unsigned(222, 10) ) ELSE
                        coeff259 WHEN ( cur_count = to_unsigned(223, 10) ) ELSE
                        coeff260 WHEN ( cur_count = to_unsigned(224, 10) ) ELSE
                        coeff261 WHEN ( cur_count = to_unsigned(225, 10) ) ELSE
                        coeff262 WHEN ( cur_count = to_unsigned(226, 10) ) ELSE
                        coeff263 WHEN ( cur_count = to_unsigned(227, 10) ) ELSE
                        coeff264 WHEN ( cur_count = to_unsigned(228, 10) ) ELSE
                        coeff265 WHEN ( cur_count = to_unsigned(229, 10) ) ELSE
                        coeff266 WHEN ( cur_count = to_unsigned(230, 10) ) ELSE
                        coeff267 WHEN ( cur_count = to_unsigned(231, 10) ) ELSE
                        coeff268 WHEN ( cur_count = to_unsigned(232, 10) ) ELSE
                        coeff269 WHEN ( cur_count = to_unsigned(233, 10) ) ELSE
                        coeff270 WHEN ( cur_count = to_unsigned(234, 10) ) ELSE
                        coeff271 WHEN ( cur_count = to_unsigned(235, 10) ) ELSE
                        coeff272 WHEN ( cur_count = to_unsigned(236, 10) ) ELSE
                        coeff273 WHEN ( cur_count = to_unsigned(237, 10) ) ELSE
                        coeff274 WHEN ( cur_count = to_unsigned(238, 10) ) ELSE
                        coeff275 WHEN ( cur_count = to_unsigned(239, 10) ) ELSE
                        coeff276 WHEN ( cur_count = to_unsigned(240, 10) ) ELSE
                        coeff277 WHEN ( cur_count = to_unsigned(241, 10) ) ELSE
                        coeff278 WHEN ( cur_count = to_unsigned(242, 10) ) ELSE
                        coeff279 WHEN ( cur_count = to_unsigned(243, 10) ) ELSE
                        coeff280 WHEN ( cur_count = to_unsigned(244, 10) ) ELSE
                        coeff281 WHEN ( cur_count = to_unsigned(245, 10) ) ELSE
                        coeff282 WHEN ( cur_count = to_unsigned(246, 10) ) ELSE
                        coeff283 WHEN ( cur_count = to_unsigned(247, 10) ) ELSE
                        coeff284 WHEN ( cur_count = to_unsigned(248, 10) ) ELSE
                        coeff285 WHEN ( cur_count = to_unsigned(249, 10) ) ELSE
                        coeff286 WHEN ( cur_count = to_unsigned(250, 10) ) ELSE
                        coeff287 WHEN ( cur_count = to_unsigned(251, 10) ) ELSE
                        coeff288 WHEN ( cur_count = to_unsigned(252, 10) ) ELSE
                        coeff289 WHEN ( cur_count = to_unsigned(253, 10) ) ELSE
                        coeff290 WHEN ( cur_count = to_unsigned(254, 10) ) ELSE
                        coeff291 WHEN ( cur_count = to_unsigned(255, 10) ) ELSE
                        coeff292 WHEN ( cur_count = to_unsigned(256, 10) ) ELSE
                        coeff293 WHEN ( cur_count = to_unsigned(257, 10) ) ELSE
                        coeff294 WHEN ( cur_count = to_unsigned(258, 10) ) ELSE
                        coeff295 WHEN ( cur_count = to_unsigned(259, 10) ) ELSE
                        coeff296 WHEN ( cur_count = to_unsigned(260, 10) ) ELSE
                        coeff297 WHEN ( cur_count = to_unsigned(261, 10) ) ELSE
                        coeff298 WHEN ( cur_count = to_unsigned(262, 10) ) ELSE
                        coeff300 WHEN ( cur_count = to_unsigned(263, 10) ) ELSE
                        coeff301 WHEN ( cur_count = to_unsigned(264, 10) ) ELSE
                        coeff302 WHEN ( cur_count = to_unsigned(265, 10) ) ELSE
                        coeff303 WHEN ( cur_count = to_unsigned(266, 10) ) ELSE
                        coeff304 WHEN ( cur_count = to_unsigned(267, 10) ) ELSE
                        coeff305 WHEN ( cur_count = to_unsigned(268, 10) ) ELSE
                        coeff306 WHEN ( cur_count = to_unsigned(269, 10) ) ELSE
                        coeff307 WHEN ( cur_count = to_unsigned(270, 10) ) ELSE
                        coeff308 WHEN ( cur_count = to_unsigned(271, 10) ) ELSE
                        coeff309 WHEN ( cur_count = to_unsigned(272, 10) ) ELSE
                        coeff310 WHEN ( cur_count = to_unsigned(273, 10) ) ELSE
                        coeff311 WHEN ( cur_count = to_unsigned(274, 10) ) ELSE
                        coeff312 WHEN ( cur_count = to_unsigned(275, 10) ) ELSE
                        coeff313 WHEN ( cur_count = to_unsigned(276, 10) ) ELSE
                        coeff314 WHEN ( cur_count = to_unsigned(277, 10) ) ELSE
                        coeff315 WHEN ( cur_count = to_unsigned(278, 10) ) ELSE
                        coeff316 WHEN ( cur_count = to_unsigned(279, 10) ) ELSE
                        coeff317 WHEN ( cur_count = to_unsigned(280, 10) ) ELSE
                        coeff318 WHEN ( cur_count = to_unsigned(281, 10) ) ELSE
                        coeff319 WHEN ( cur_count = to_unsigned(282, 10) ) ELSE
                        coeff320 WHEN ( cur_count = to_unsigned(283, 10) ) ELSE
                        coeff321 WHEN ( cur_count = to_unsigned(284, 10) ) ELSE
                        coeff322 WHEN ( cur_count = to_unsigned(285, 10) ) ELSE
                        coeff323 WHEN ( cur_count = to_unsigned(286, 10) ) ELSE
                        coeff324 WHEN ( cur_count = to_unsigned(287, 10) ) ELSE
                        coeff325 WHEN ( cur_count = to_unsigned(288, 10) ) ELSE
                        coeff326 WHEN ( cur_count = to_unsigned(289, 10) ) ELSE
                        coeff327 WHEN ( cur_count = to_unsigned(290, 10) ) ELSE
                        coeff328 WHEN ( cur_count = to_unsigned(291, 10) ) ELSE
                        coeff329 WHEN ( cur_count = to_unsigned(292, 10) ) ELSE
                        coeff330 WHEN ( cur_count = to_unsigned(293, 10) ) ELSE
                        coeff331 WHEN ( cur_count = to_unsigned(294, 10) ) ELSE
                        coeff332 WHEN ( cur_count = to_unsigned(295, 10) ) ELSE
                        coeff333 WHEN ( cur_count = to_unsigned(296, 10) ) ELSE
                        coeff334 WHEN ( cur_count = to_unsigned(297, 10) ) ELSE
                        coeff335 WHEN ( cur_count = to_unsigned(298, 10) ) ELSE
                        coeff336 WHEN ( cur_count = to_unsigned(299, 10) ) ELSE
                        coeff337 WHEN ( cur_count = to_unsigned(300, 10) ) ELSE
                        coeff338 WHEN ( cur_count = to_unsigned(301, 10) ) ELSE
                        coeff339 WHEN ( cur_count = to_unsigned(302, 10) ) ELSE
                        coeff340 WHEN ( cur_count = to_unsigned(303, 10) ) ELSE
                        coeff341 WHEN ( cur_count = to_unsigned(304, 10) ) ELSE
                        coeff342 WHEN ( cur_count = to_unsigned(305, 10) ) ELSE
                        coeff343 WHEN ( cur_count = to_unsigned(306, 10) ) ELSE
                        coeff344 WHEN ( cur_count = to_unsigned(307, 10) ) ELSE
                        coeff345 WHEN ( cur_count = to_unsigned(308, 10) ) ELSE
                        coeff346 WHEN ( cur_count = to_unsigned(309, 10) ) ELSE
                        coeff347 WHEN ( cur_count = to_unsigned(310, 10) ) ELSE
                        coeff348 WHEN ( cur_count = to_unsigned(311, 10) ) ELSE
                        coeff349 WHEN ( cur_count = to_unsigned(312, 10) ) ELSE
                        coeff350 WHEN ( cur_count = to_unsigned(313, 10) ) ELSE
                        coeff351 WHEN ( cur_count = to_unsigned(314, 10) ) ELSE
                        coeff352 WHEN ( cur_count = to_unsigned(315, 10) ) ELSE
                        coeff353 WHEN ( cur_count = to_unsigned(316, 10) ) ELSE
                        coeff354 WHEN ( cur_count = to_unsigned(317, 10) ) ELSE
                        coeff355 WHEN ( cur_count = to_unsigned(318, 10) ) ELSE
                        coeff356 WHEN ( cur_count = to_unsigned(319, 10) ) ELSE
                        coeff357 WHEN ( cur_count = to_unsigned(320, 10) ) ELSE
                        coeff358 WHEN ( cur_count = to_unsigned(321, 10) ) ELSE
                        coeff359 WHEN ( cur_count = to_unsigned(322, 10) ) ELSE
                        coeff360 WHEN ( cur_count = to_unsigned(323, 10) ) ELSE
                        coeff361 WHEN ( cur_count = to_unsigned(324, 10) ) ELSE
                        coeff362 WHEN ( cur_count = to_unsigned(325, 10) ) ELSE
                        coeff363 WHEN ( cur_count = to_unsigned(326, 10) ) ELSE
                        coeff364 WHEN ( cur_count = to_unsigned(327, 10) ) ELSE
                        coeff365 WHEN ( cur_count = to_unsigned(328, 10) ) ELSE
                        coeff366 WHEN ( cur_count = to_unsigned(329, 10) ) ELSE
                        coeff367 WHEN ( cur_count = to_unsigned(330, 10) ) ELSE
                        coeff368 WHEN ( cur_count = to_unsigned(331, 10) ) ELSE
                        coeff369 WHEN ( cur_count = to_unsigned(332, 10) ) ELSE
                        coeff370 WHEN ( cur_count = to_unsigned(333, 10) ) ELSE
                        coeff371 WHEN ( cur_count = to_unsigned(334, 10) ) ELSE
                        coeff372 WHEN ( cur_count = to_unsigned(335, 10) ) ELSE
                        coeff373 WHEN ( cur_count = to_unsigned(336, 10) ) ELSE
                        coeff374 WHEN ( cur_count = to_unsigned(337, 10) ) ELSE
                        coeff375 WHEN ( cur_count = to_unsigned(338, 10) ) ELSE
                        coeff376 WHEN ( cur_count = to_unsigned(339, 10) ) ELSE
                        coeff377 WHEN ( cur_count = to_unsigned(340, 10) ) ELSE
                        coeff378 WHEN ( cur_count = to_unsigned(341, 10) ) ELSE
                        coeff379 WHEN ( cur_count = to_unsigned(342, 10) ) ELSE
                        coeff380 WHEN ( cur_count = to_unsigned(343, 10) ) ELSE
                        coeff381 WHEN ( cur_count = to_unsigned(344, 10) ) ELSE
                        coeff382 WHEN ( cur_count = to_unsigned(345, 10) ) ELSE
                        coeff383 WHEN ( cur_count = to_unsigned(346, 10) ) ELSE
                        coeff384 WHEN ( cur_count = to_unsigned(347, 10) ) ELSE
                        coeff385 WHEN ( cur_count = to_unsigned(348, 10) ) ELSE
                        coeff386 WHEN ( cur_count = to_unsigned(349, 10) ) ELSE
                        coeff387 WHEN ( cur_count = to_unsigned(350, 10) ) ELSE
                        coeff388 WHEN ( cur_count = to_unsigned(351, 10) ) ELSE
                        coeff389 WHEN ( cur_count = to_unsigned(352, 10) ) ELSE
                        coeff390 WHEN ( cur_count = to_unsigned(353, 10) ) ELSE
                        coeff391 WHEN ( cur_count = to_unsigned(354, 10) ) ELSE
                        coeff392 WHEN ( cur_count = to_unsigned(355, 10) ) ELSE
                        coeff393 WHEN ( cur_count = to_unsigned(356, 10) ) ELSE
                        coeff394 WHEN ( cur_count = to_unsigned(357, 10) ) ELSE
                        coeff395 WHEN ( cur_count = to_unsigned(358, 10) ) ELSE
                        coeff397 WHEN ( cur_count = to_unsigned(359, 10) ) ELSE
                        coeff398 WHEN ( cur_count = to_unsigned(360, 10) ) ELSE
                        coeff399 WHEN ( cur_count = to_unsigned(361, 10) ) ELSE
                        coeff400 WHEN ( cur_count = to_unsigned(362, 10) ) ELSE
                        coeff401 WHEN ( cur_count = to_unsigned(363, 10) ) ELSE
                        coeff402 WHEN ( cur_count = to_unsigned(364, 10) ) ELSE
                        coeff403 WHEN ( cur_count = to_unsigned(365, 10) ) ELSE
                        coeff404 WHEN ( cur_count = to_unsigned(366, 10) ) ELSE
                        coeff405 WHEN ( cur_count = to_unsigned(367, 10) ) ELSE
                        coeff406 WHEN ( cur_count = to_unsigned(368, 10) ) ELSE
                        coeff407 WHEN ( cur_count = to_unsigned(369, 10) ) ELSE
                        coeff408 WHEN ( cur_count = to_unsigned(370, 10) ) ELSE
                        coeff409 WHEN ( cur_count = to_unsigned(371, 10) ) ELSE
                        coeff410 WHEN ( cur_count = to_unsigned(372, 10) ) ELSE
                        coeff411 WHEN ( cur_count = to_unsigned(373, 10) ) ELSE
                        coeff412 WHEN ( cur_count = to_unsigned(374, 10) ) ELSE
                        coeff413 WHEN ( cur_count = to_unsigned(375, 10) ) ELSE
                        coeff414 WHEN ( cur_count = to_unsigned(376, 10) ) ELSE
                        coeff415 WHEN ( cur_count = to_unsigned(377, 10) ) ELSE
                        coeff416 WHEN ( cur_count = to_unsigned(378, 10) ) ELSE
                        coeff417 WHEN ( cur_count = to_unsigned(379, 10) ) ELSE
                        coeff418 WHEN ( cur_count = to_unsigned(380, 10) ) ELSE
                        coeff419 WHEN ( cur_count = to_unsigned(381, 10) ) ELSE
                        coeff420 WHEN ( cur_count = to_unsigned(382, 10) ) ELSE
                        coeff421 WHEN ( cur_count = to_unsigned(383, 10) ) ELSE
                        coeff422 WHEN ( cur_count = to_unsigned(384, 10) ) ELSE
                        coeff423 WHEN ( cur_count = to_unsigned(385, 10) ) ELSE
                        coeff424 WHEN ( cur_count = to_unsigned(386, 10) ) ELSE
                        coeff425 WHEN ( cur_count = to_unsigned(387, 10) ) ELSE
                        coeff426 WHEN ( cur_count = to_unsigned(388, 10) ) ELSE
                        coeff427 WHEN ( cur_count = to_unsigned(389, 10) ) ELSE
                        coeff428 WHEN ( cur_count = to_unsigned(390, 10) ) ELSE
                        coeff429 WHEN ( cur_count = to_unsigned(391, 10) ) ELSE
                        coeff430 WHEN ( cur_count = to_unsigned(392, 10) ) ELSE
                        coeff431 WHEN ( cur_count = to_unsigned(393, 10) ) ELSE
                        coeff432 WHEN ( cur_count = to_unsigned(394, 10) ) ELSE
                        coeff433 WHEN ( cur_count = to_unsigned(395, 10) ) ELSE
                        coeff434 WHEN ( cur_count = to_unsigned(396, 10) ) ELSE
                        coeff435 WHEN ( cur_count = to_unsigned(397, 10) ) ELSE
                        coeff436 WHEN ( cur_count = to_unsigned(398, 10) ) ELSE
                        coeff437 WHEN ( cur_count = to_unsigned(399, 10) ) ELSE
                        coeff438 WHEN ( cur_count = to_unsigned(400, 10) ) ELSE
                        coeff439 WHEN ( cur_count = to_unsigned(401, 10) ) ELSE
                        coeff440 WHEN ( cur_count = to_unsigned(402, 10) ) ELSE
                        coeff441 WHEN ( cur_count = to_unsigned(403, 10) ) ELSE
                        coeff442 WHEN ( cur_count = to_unsigned(404, 10) ) ELSE
                        coeff443 WHEN ( cur_count = to_unsigned(405, 10) ) ELSE
                        coeff445 WHEN ( cur_count = to_unsigned(406, 10) ) ELSE
                        coeff446 WHEN ( cur_count = to_unsigned(407, 10) ) ELSE
                        coeff447 WHEN ( cur_count = to_unsigned(408, 10) ) ELSE
                        coeff448 WHEN ( cur_count = to_unsigned(409, 10) ) ELSE
                        coeff449 WHEN ( cur_count = to_unsigned(410, 10) ) ELSE
                        coeff450 WHEN ( cur_count = to_unsigned(411, 10) ) ELSE
                        coeff451 WHEN ( cur_count = to_unsigned(412, 10) ) ELSE
                        coeff452 WHEN ( cur_count = to_unsigned(413, 10) ) ELSE
                        coeff453 WHEN ( cur_count = to_unsigned(414, 10) ) ELSE
                        coeff454 WHEN ( cur_count = to_unsigned(415, 10) ) ELSE
                        coeff455 WHEN ( cur_count = to_unsigned(416, 10) ) ELSE
                        coeff456 WHEN ( cur_count = to_unsigned(417, 10) ) ELSE
                        coeff457 WHEN ( cur_count = to_unsigned(418, 10) ) ELSE
                        coeff458 WHEN ( cur_count = to_unsigned(419, 10) ) ELSE
                        coeff459 WHEN ( cur_count = to_unsigned(420, 10) ) ELSE
                        coeff460 WHEN ( cur_count = to_unsigned(421, 10) ) ELSE
                        coeff461 WHEN ( cur_count = to_unsigned(422, 10) ) ELSE
                        coeff462 WHEN ( cur_count = to_unsigned(423, 10) ) ELSE
                        coeff463 WHEN ( cur_count = to_unsigned(424, 10) ) ELSE
                        coeff464 WHEN ( cur_count = to_unsigned(425, 10) ) ELSE
                        coeff465 WHEN ( cur_count = to_unsigned(426, 10) ) ELSE
                        coeff466 WHEN ( cur_count = to_unsigned(427, 10) ) ELSE
                        coeff467 WHEN ( cur_count = to_unsigned(428, 10) ) ELSE
                        coeff468 WHEN ( cur_count = to_unsigned(429, 10) ) ELSE
                        coeff469 WHEN ( cur_count = to_unsigned(430, 10) ) ELSE
                        coeff470 WHEN ( cur_count = to_unsigned(431, 10) ) ELSE
                        coeff471 WHEN ( cur_count = to_unsigned(432, 10) ) ELSE
                        coeff472 WHEN ( cur_count = to_unsigned(433, 10) ) ELSE
                        coeff473 WHEN ( cur_count = to_unsigned(434, 10) ) ELSE
                        coeff474 WHEN ( cur_count = to_unsigned(435, 10) ) ELSE
                        coeff475 WHEN ( cur_count = to_unsigned(436, 10) ) ELSE
                        coeff476 WHEN ( cur_count = to_unsigned(437, 10) ) ELSE
                        coeff477 WHEN ( cur_count = to_unsigned(438, 10) ) ELSE
                        coeff478 WHEN ( cur_count = to_unsigned(439, 10) ) ELSE
                        coeff479 WHEN ( cur_count = to_unsigned(440, 10) ) ELSE
                        coeff480 WHEN ( cur_count = to_unsigned(441, 10) ) ELSE
                        coeff481 WHEN ( cur_count = to_unsigned(442, 10) ) ELSE
                        coeff482 WHEN ( cur_count = to_unsigned(443, 10) ) ELSE
                        coeff483 WHEN ( cur_count = to_unsigned(444, 10) ) ELSE
                        coeff484 WHEN ( cur_count = to_unsigned(445, 10) ) ELSE
                        coeff485 WHEN ( cur_count = to_unsigned(446, 10) ) ELSE
                        coeff486 WHEN ( cur_count = to_unsigned(447, 10) ) ELSE
                        coeff487 WHEN ( cur_count = to_unsigned(448, 10) ) ELSE
                        coeff488 WHEN ( cur_count = to_unsigned(449, 10) ) ELSE
                        coeff489 WHEN ( cur_count = to_unsigned(450, 10) ) ELSE
                        coeff490 WHEN ( cur_count = to_unsigned(451, 10) ) ELSE
                        coeff491 WHEN ( cur_count = to_unsigned(452, 10) ) ELSE
                        coeff494 WHEN ( cur_count = to_unsigned(453, 10) ) ELSE
                        coeff495 WHEN ( cur_count = to_unsigned(454, 10) ) ELSE
                        coeff496 WHEN ( cur_count = to_unsigned(455, 10) ) ELSE
                        coeff497 WHEN ( cur_count = to_unsigned(456, 10) ) ELSE
                        coeff498 WHEN ( cur_count = to_unsigned(457, 10) ) ELSE
                        coeff499 WHEN ( cur_count = to_unsigned(458, 10) ) ELSE
                        coeff500 WHEN ( cur_count = to_unsigned(459, 10) ) ELSE
                        coeff501 WHEN ( cur_count = to_unsigned(460, 10) ) ELSE
                        coeff502 WHEN ( cur_count = to_unsigned(461, 10) ) ELSE
                        coeff503 WHEN ( cur_count = to_unsigned(462, 10) ) ELSE
                        coeff504 WHEN ( cur_count = to_unsigned(463, 10) ) ELSE
                        coeff505 WHEN ( cur_count = to_unsigned(464, 10) ) ELSE
                        coeff506 WHEN ( cur_count = to_unsigned(465, 10) ) ELSE
                        coeff507 WHEN ( cur_count = to_unsigned(466, 10) ) ELSE
                        coeff508 WHEN ( cur_count = to_unsigned(467, 10) ) ELSE
                        coeff509 WHEN ( cur_count = to_unsigned(468, 10) ) ELSE
                        coeff510 WHEN ( cur_count = to_unsigned(469, 10) ) ELSE
                        coeff511 WHEN ( cur_count = to_unsigned(470, 10) ) ELSE
                        coeff512 WHEN ( cur_count = to_unsigned(471, 10) ) ELSE
                        coeff513 WHEN ( cur_count = to_unsigned(472, 10) ) ELSE
                        coeff514 WHEN ( cur_count = to_unsigned(473, 10) ) ELSE
                        coeff515 WHEN ( cur_count = to_unsigned(474, 10) ) ELSE
                        coeff516 WHEN ( cur_count = to_unsigned(475, 10) ) ELSE
                        coeff517 WHEN ( cur_count = to_unsigned(476, 10) ) ELSE
                        coeff518 WHEN ( cur_count = to_unsigned(477, 10) ) ELSE
                        coeff519 WHEN ( cur_count = to_unsigned(478, 10) ) ELSE
                        coeff520 WHEN ( cur_count = to_unsigned(479, 10) ) ELSE
                        coeff521 WHEN ( cur_count = to_unsigned(480, 10) ) ELSE
                        coeff522 WHEN ( cur_count = to_unsigned(481, 10) ) ELSE
                        coeff523 WHEN ( cur_count = to_unsigned(482, 10) ) ELSE
                        coeff524 WHEN ( cur_count = to_unsigned(483, 10) ) ELSE
                        coeff525 WHEN ( cur_count = to_unsigned(484, 10) ) ELSE
                        coeff526 WHEN ( cur_count = to_unsigned(485, 10) ) ELSE
                        coeff527 WHEN ( cur_count = to_unsigned(486, 10) ) ELSE
                        coeff528 WHEN ( cur_count = to_unsigned(487, 10) ) ELSE
                        coeff529 WHEN ( cur_count = to_unsigned(488, 10) ) ELSE
                        coeff530 WHEN ( cur_count = to_unsigned(489, 10) ) ELSE
                        coeff531 WHEN ( cur_count = to_unsigned(490, 10) ) ELSE
                        coeff532 WHEN ( cur_count = to_unsigned(491, 10) ) ELSE
                        coeff533 WHEN ( cur_count = to_unsigned(492, 10) ) ELSE
                        coeff534 WHEN ( cur_count = to_unsigned(493, 10) ) ELSE
                        coeff535 WHEN ( cur_count = to_unsigned(494, 10) ) ELSE
                        coeff536 WHEN ( cur_count = to_unsigned(495, 10) ) ELSE
                        coeff537 WHEN ( cur_count = to_unsigned(496, 10) ) ELSE
                        coeff538 WHEN ( cur_count = to_unsigned(497, 10) ) ELSE
                        coeff543 WHEN ( cur_count = to_unsigned(498, 10) ) ELSE
                        coeff544 WHEN ( cur_count = to_unsigned(499, 10) ) ELSE
                        coeff545 WHEN ( cur_count = to_unsigned(500, 10) ) ELSE
                        coeff546 WHEN ( cur_count = to_unsigned(501, 10) ) ELSE
                        coeff547 WHEN ( cur_count = to_unsigned(502, 10) ) ELSE
                        coeff548 WHEN ( cur_count = to_unsigned(503, 10) ) ELSE
                        coeff549 WHEN ( cur_count = to_unsigned(504, 10) ) ELSE
                        coeff550 WHEN ( cur_count = to_unsigned(505, 10) ) ELSE
                        coeff551 WHEN ( cur_count = to_unsigned(506, 10) ) ELSE
                        coeff552 WHEN ( cur_count = to_unsigned(507, 10) ) ELSE
                        coeff553 WHEN ( cur_count = to_unsigned(508, 10) ) ELSE
                        coeff554 WHEN ( cur_count = to_unsigned(509, 10) ) ELSE
                        coeff555 WHEN ( cur_count = to_unsigned(510, 10) ) ELSE
                        coeff556 WHEN ( cur_count = to_unsigned(511, 10) ) ELSE
                        coeff557 WHEN ( cur_count = to_unsigned(512, 10) ) ELSE
                        coeff558 WHEN ( cur_count = to_unsigned(513, 10) ) ELSE
                        coeff559 WHEN ( cur_count = to_unsigned(514, 10) ) ELSE
                        coeff560 WHEN ( cur_count = to_unsigned(515, 10) ) ELSE
                        coeff561 WHEN ( cur_count = to_unsigned(516, 10) ) ELSE
                        coeff562 WHEN ( cur_count = to_unsigned(517, 10) ) ELSE
                        coeff563 WHEN ( cur_count = to_unsigned(518, 10) ) ELSE
                        coeff564 WHEN ( cur_count = to_unsigned(519, 10) ) ELSE
                        coeff565 WHEN ( cur_count = to_unsigned(520, 10) ) ELSE
                        coeff566 WHEN ( cur_count = to_unsigned(521, 10) ) ELSE
                        coeff567 WHEN ( cur_count = to_unsigned(522, 10) ) ELSE
                        coeff568 WHEN ( cur_count = to_unsigned(523, 10) ) ELSE
                        coeff569 WHEN ( cur_count = to_unsigned(524, 10) ) ELSE
                        coeff570 WHEN ( cur_count = to_unsigned(525, 10) ) ELSE
                        coeff571 WHEN ( cur_count = to_unsigned(526, 10) ) ELSE
                        coeff572 WHEN ( cur_count = to_unsigned(527, 10) ) ELSE
                        coeff573 WHEN ( cur_count = to_unsigned(528, 10) ) ELSE
                        coeff574 WHEN ( cur_count = to_unsigned(529, 10) ) ELSE
                        coeff575 WHEN ( cur_count = to_unsigned(530, 10) ) ELSE
                        coeff576 WHEN ( cur_count = to_unsigned(531, 10) ) ELSE
                        coeff577 WHEN ( cur_count = to_unsigned(532, 10) ) ELSE
                        coeff578 WHEN ( cur_count = to_unsigned(533, 10) ) ELSE
                        coeff579 WHEN ( cur_count = to_unsigned(534, 10) ) ELSE
                        coeff580 WHEN ( cur_count = to_unsigned(535, 10) ) ELSE
                        coeff581 WHEN ( cur_count = to_unsigned(536, 10) ) ELSE
                        coeff582 WHEN ( cur_count = to_unsigned(537, 10) ) ELSE
                        coeff583 WHEN ( cur_count = to_unsigned(538, 10) ) ELSE
                        coeff584 WHEN ( cur_count = to_unsigned(539, 10) ) ELSE
                        coeff592 WHEN ( cur_count = to_unsigned(540, 10) ) ELSE
                        coeff593 WHEN ( cur_count = to_unsigned(541, 10) ) ELSE
                        coeff594 WHEN ( cur_count = to_unsigned(542, 10) ) ELSE
                        coeff595 WHEN ( cur_count = to_unsigned(543, 10) ) ELSE
                        coeff596 WHEN ( cur_count = to_unsigned(544, 10) ) ELSE
                        coeff597 WHEN ( cur_count = to_unsigned(545, 10) ) ELSE
                        coeff598 WHEN ( cur_count = to_unsigned(546, 10) ) ELSE
                        coeff599 WHEN ( cur_count = to_unsigned(547, 10) ) ELSE
                        coeff600 WHEN ( cur_count = to_unsigned(548, 10) ) ELSE
                        coeff601 WHEN ( cur_count = to_unsigned(549, 10) ) ELSE
                        coeff602 WHEN ( cur_count = to_unsigned(550, 10) ) ELSE
                        coeff603 WHEN ( cur_count = to_unsigned(551, 10) ) ELSE
                        coeff604 WHEN ( cur_count = to_unsigned(552, 10) ) ELSE
                        coeff605 WHEN ( cur_count = to_unsigned(553, 10) ) ELSE
                        coeff606 WHEN ( cur_count = to_unsigned(554, 10) ) ELSE
                        coeff607 WHEN ( cur_count = to_unsigned(555, 10) ) ELSE
                        coeff608 WHEN ( cur_count = to_unsigned(556, 10) ) ELSE
                        coeff609 WHEN ( cur_count = to_unsigned(557, 10) ) ELSE
                        coeff610 WHEN ( cur_count = to_unsigned(558, 10) ) ELSE
                        coeff611 WHEN ( cur_count = to_unsigned(559, 10) ) ELSE
                        coeff612 WHEN ( cur_count = to_unsigned(560, 10) ) ELSE
                        coeff613 WHEN ( cur_count = to_unsigned(561, 10) ) ELSE
                        coeff614 WHEN ( cur_count = to_unsigned(562, 10) ) ELSE
                        coeff615 WHEN ( cur_count = to_unsigned(563, 10) ) ELSE
                        coeff616 WHEN ( cur_count = to_unsigned(564, 10) ) ELSE
                        coeff617 WHEN ( cur_count = to_unsigned(565, 10) ) ELSE
                        coeff618 WHEN ( cur_count = to_unsigned(566, 10) ) ELSE
                        coeff619 WHEN ( cur_count = to_unsigned(567, 10) ) ELSE
                        coeff620 WHEN ( cur_count = to_unsigned(568, 10) ) ELSE
                        coeff621 WHEN ( cur_count = to_unsigned(569, 10) ) ELSE
                        coeff622 WHEN ( cur_count = to_unsigned(570, 10) ) ELSE
                        coeff623 WHEN ( cur_count = to_unsigned(571, 10) ) ELSE
                        coeff624 WHEN ( cur_count = to_unsigned(572, 10) ) ELSE
                        coeff625 WHEN ( cur_count = to_unsigned(573, 10) ) ELSE
                        coeff626 WHEN ( cur_count = to_unsigned(574, 10) ) ELSE
                        coeff627 WHEN ( cur_count = to_unsigned(575, 10) ) ELSE
                        coeff628 WHEN ( cur_count = to_unsigned(576, 10) ) ELSE
                        coeff629 WHEN ( cur_count = to_unsigned(577, 10) ) ELSE
                        coeff643 WHEN ( cur_count = to_unsigned(578, 10) ) ELSE
                        coeff644 WHEN ( cur_count = to_unsigned(579, 10) ) ELSE
                        coeff645 WHEN ( cur_count = to_unsigned(580, 10) ) ELSE
                        coeff646 WHEN ( cur_count = to_unsigned(581, 10) ) ELSE
                        coeff647 WHEN ( cur_count = to_unsigned(582, 10) ) ELSE
                        coeff648 WHEN ( cur_count = to_unsigned(583, 10) ) ELSE
                        coeff649 WHEN ( cur_count = to_unsigned(584, 10) ) ELSE
                        coeff650 WHEN ( cur_count = to_unsigned(585, 10) ) ELSE
                        coeff651 WHEN ( cur_count = to_unsigned(586, 10) ) ELSE
                        coeff652 WHEN ( cur_count = to_unsigned(587, 10) ) ELSE
                        coeff653 WHEN ( cur_count = to_unsigned(588, 10) ) ELSE
                        coeff654 WHEN ( cur_count = to_unsigned(589, 10) ) ELSE
                        coeff655 WHEN ( cur_count = to_unsigned(590, 10) ) ELSE
                        coeff656 WHEN ( cur_count = to_unsigned(591, 10) ) ELSE
                        coeff657 WHEN ( cur_count = to_unsigned(592, 10) ) ELSE
                        coeff658 WHEN ( cur_count = to_unsigned(593, 10) ) ELSE
                        coeff659 WHEN ( cur_count = to_unsigned(594, 10) ) ELSE
                        coeff660 WHEN ( cur_count = to_unsigned(595, 10) ) ELSE
                        coeff661 WHEN ( cur_count = to_unsigned(596, 10) ) ELSE
                        coeff662 WHEN ( cur_count = to_unsigned(597, 10) ) ELSE
                        coeff663 WHEN ( cur_count = to_unsigned(598, 10) ) ELSE
                        coeff664 WHEN ( cur_count = to_unsigned(599, 10) ) ELSE
                        coeff665 WHEN ( cur_count = to_unsigned(600, 10) ) ELSE
                        coeff666 WHEN ( cur_count = to_unsigned(601, 10) ) ELSE
                        coeff667 WHEN ( cur_count = to_unsigned(602, 10) ) ELSE
                        coeff668 WHEN ( cur_count = to_unsigned(603, 10) ) ELSE
                        coeff669 WHEN ( cur_count = to_unsigned(604, 10) ) ELSE
                        coeff670 WHEN ( cur_count = to_unsigned(605, 10) ) ELSE
                        coeff671 WHEN ( cur_count = to_unsigned(606, 10) ) ELSE
                        coeff672 WHEN ( cur_count = to_unsigned(607, 10) ) ELSE
                        coeff673 WHEN ( cur_count = to_unsigned(608, 10) ) ELSE
                        coeff674 WHEN ( cur_count = to_unsigned(609, 10) ) ELSE
                        coeff675 WHEN ( cur_count = to_unsigned(610, 10) ) ELSE
                        coeff676 WHEN ( cur_count = to_unsigned(611, 10) ) ELSE
                        coeff677 WHEN ( cur_count = to_unsigned(612, 10) ) ELSE
                        coeff686 WHEN ( cur_count = to_unsigned(613, 10) ) ELSE
                        coeff687 WHEN ( cur_count = to_unsigned(614, 10) ) ELSE
                        coeff688 WHEN ( cur_count = to_unsigned(615, 10) ) ELSE
                        coeff689 WHEN ( cur_count = to_unsigned(616, 10) ) ELSE
                        coeff690 WHEN ( cur_count = to_unsigned(617, 10) ) ELSE
                        coeff691 WHEN ( cur_count = to_unsigned(618, 10) ) ELSE
                        coeff692 WHEN ( cur_count = to_unsigned(619, 10) ) ELSE
                        coeff693 WHEN ( cur_count = to_unsigned(620, 10) ) ELSE
                        coeff694;
  mul_temp <= inputmux_1 * product_1_mux;
  product_1 <= mul_temp(38 DOWNTO 0);

  prod_typeconvert_1 <= resize(product_1, 45);

  add_temp <= resize(prod_typeconvert_1, 46) + resize(acc_out_1, 46);
  acc_sum_1 <= add_temp(44 DOWNTO 0);

  acc_in_1 <= prod_typeconvert_1 WHEN ( phase_0 = '1' ) ELSE
                   acc_sum_1;

  Acc_reg_1_process : PROCESS (I_CLK, I_RST)
  BEGIN
    IF I_RST = '1' THEN
      acc_out_1 <= (OTHERS => '0');
    ELSIF rising_edge(I_CLK) THEN
      acc_out_1 <= acc_in_1;
    END IF;
  END PROCESS Acc_reg_1_process;

  Finalsum_reg_process : PROCESS (I_CLK, I_RST)
  BEGIN
    IF I_RST = '1' THEN
      acc_final <= (OTHERS => '0');
    ELSIF rising_edge(I_CLK) THEN
      IF phase_0 = '1' THEN
        acc_final <= acc_out_1;
      END IF;
    END IF;
  END PROCESS Finalsum_reg_process;

  output_typeconvert <= acc_final;

  Output_Register_process : PROCESS (I_CLK, I_RST)
  BEGIN
    IF I_RST = '1' THEN
      output_register <= (OTHERS => '0');
    ELSIF rising_edge(I_CLK) THEN
      IF phase_0 = '1' THEN
        output_register <= output_typeconvert;
      END IF;
    END IF;
  END PROCESS Output_Register_process;

  -- Assignment Statements
  O_FILTER <= std_logic_vector(output_register);
END architecture rtl;