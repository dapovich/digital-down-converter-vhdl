------------------------------------------------------------------
--  File        : dpROM12.vhd
--  Description : Direct Digital Synthesis top level
------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity hf_generator is
  port (
    I_CLK : in std_logic;
    I_RST : in std_logic;
    I_PHASEINC : in std_logic_vector(31 downto 0);
    O_SINE : out std_logic_vector(15 downto 0)
  );
end entity hf_generator;

architecture rtl of hf_generator is

  -- Initialize sine Look-up table ROM component
  component dpROM12 is
  port (
    I_CLK    : in std_logic;
    I_ADDR_A : in std_logic_vector(9 downto 0);
    I_ADDR_B : in std_logic_vector(9 downto 0);
    O_DATA_A : out std_logic_vector(15 downto 0);
    O_DATA_B : out std_logic_vector(15 downto 0)
  );
  end component dpROM12;

  -- Internal signals
  signal tuningWord_reg : std_logic_vector(31 downto 0) := (others => '0');
  signal phaseAccum : unsigned(31 downto 0) := (others => '0');
  signal ditherWord : unsigned(31 downto 0) := (others => '0');
  signal lfsrWord   : unsigned(31 downto 0) := x"00000001";
  signal addrDelay  : std_logic_vector(31 downto 30) := "00";

  signal sin : std_logic_vector(15 downto 0);
  signal romAddr_sin : std_logic_vector(9 downto 0);
  signal sin_invert : std_logic_vector(15 downto 0);
  signal sin_2s_comp : unsigned(15 downto 0);
  signal sinwave : std_logic_vector(15 downto 0);

  signal empty_16 : std_logic_vector(15 downto 0);
  signal empty_10 : std_logic_vector(9 downto 0) := (others => '0');
  signal cos_invert : std_logic_vector(15 downto 0);
  signal cos_2s_comp : unsigned(15 downto 0);
  signal coswave : std_logic_vector(15 downto 0) := x"7FFF";

begin

  ----------------------------------------------------------------------
  -- Instantiate Sine Look-up table
  -- @Info: sine Look-up table is a quarter-wave table to reduce memory
  -- requirements. The ROM is dual-port to allow both sin & cos to be
  -- generated
  ----------------------------------------------------------------------
  UUT : dpROM12
    port map (
      I_CLK => I_CLK,
      I_ADDR_A => romAddr_sin,
      O_DATA_A => sin,
      I_ADDR_B => empty_10,
      O_DATA_B => empty_16
  );

  ------------------------------------------
  -- 32bit Phase Accumulator
  -- For a 12bit address LUT, the phase
  -- accumulator has 20 fractional bits (19:0)
  ------------------------------------------

  -- @Task: Load tuning word to internal register
  process (I_CLK) is
  begin
    if (rising_edge(I_CLK)) then
      if (I_RST = '1') then
        tuningWord_reg <= (others => '0');
      else
        tuningWord_reg <= I_PHASEINC;
      end if;
    end if;
  end process;

  -- @Task: Phase Accumulator process
  process (I_CLK) is
  begin
    if (rising_edge(I_CLK)) then
      if (I_RST = '1') then
        phaseAccum <= (others => '0');
      else
        phaseAccum <= phaseAccum + unsigned(tuningWord_reg);
      end if;
    end if;
  end process;
  ------------------------------------------
  -- ./32bit Phase Accumulator
  ------------------------------------------

  ------------------------------------------------------------------
  -- Phase dithering
  -- A pseudo-random value is generated by a maximal length
  -- Linear Feedback Shift Register which is added to the fractional
  -- bits of the phase accumulator
  ------------------------------------------------------------------

  -- maximal length 20 bit LFSR
  process (I_CLK)
  begin
    if (rising_edge(I_CLK)) then
      lfsrWord(19 downto 1) <= lfsrWord(18 downto 0);
      lfsrWord(0) <= lfsrWord(2) xor lfsrWord(19);
    end if;
  end process;

  -- add LFSR to phase accumulator output
  process (I_CLK)
  begin
    if (rising_edge(I_CLK)) then
      if (I_RST = '1') then
        ditherWord <= (others => '0');
      else
        ditherWord <= phaseAccum + lfsrWord;
      end if;
    end if;
  end process;

  process (I_CLK)
  begin
    if (rising_edge(I_CLK)) then
      if (I_RST = '1') then
        addrDelay <= "00";
      else
        addrDelay <= std_logic_vector(phaseAccum(31 downto 30));
      end if;
    end if;
  end process;
  ------------------------------------------
  -- ./Phase dithering
  ------------------------------------------

  ------------------------------------------------------------------
  -- Sine table address
  -- The quadrant of the sine wave is selected by the 2 MS bits
  -- of the dithered phase accumulator.

  -- ditherWord (31:30)         quadrant
  ---------------------------------------------
  --       00                 0     -> pi/2
  --       01                 pi/2  -> pi
  --       10                 pi    -> 3pi/2
  --       10                 3pi/2 -> 2pi
  ------------------------------------------------------------------
  process (ditherWord)
  begin
    for i in 0 to 9 loop
      romAddr_sin(i) <= ditherWord(i+20) xor ditherWord(30);
    end loop;
  end process;
  ------------------------------------------
  -- ./Sine table address
  ------------------------------------------


  ------------------------------------------
  -- 2s Complement of sine output
  ------------------------------------------
  sin_invert <= not(sin);
  sin_2s_comp <= unsigned(sin_invert) + 1;

  process (I_CLK)
  begin
    if (rising_edge(I_CLK)) then
      if (I_RST = '1') then
        sinwave <= (others => '0');
      elsif (addrDelay(31) = '1') then
        sinwave <= std_logic_vector(sin_2s_comp);
      else
        sinwave <= sin;
      end if;
    end if;
  end process;

  O_SINE <= sinwave;
  ------------------------------------------
  -- ./2s Complement of sine output
  ------------------------------------------

end architecture rtl;

------------------------------------------------------------------
--  End of File: dpROM12.vhd
------------------------------------------------------------------

